 `include "global.sv"
`include "timescale.sv"

module sign_mnist(
	input			clk,
	input			rstn,
	input			en,
	input			go,
	
	output	reg			ready,
	output			[`WD:0]	q_data
	);
	reg	[`WD:0]		dt;
	
	reg	[1:0]		din;
	reg			push;
	
	reg	[1:0]		count;
	
	reg	[10:0]		cnt;
	reg			cnt_en;
	wire			cnt_max = cnt == 10'd783;
	wire			end_cnt_en = cnt_max;

	always @(posedge clk, negedge rstn) begin
		if(rstn == 0) begin
			din	<=	2'd0;
			push	<=	1'b0;
		end
		else begin
			if(en == 1) begin
				din[0]	<=	go;
				din[1]	<=	din[0];
				if(din[0] == 1 && din[1] == 0) begin
					push	<=	1'b1;
				end
				else begin
					push	<=	1'b0;
				end
			end
			else begin
				din	<=	2'b0;
				push	<=	1'b0;
			end
		end
	end

	always @(posedge clk, negedge rstn) begin
		if (rstn == 0) begin
			count	<=	2'd3;
		end
		else begin
			if(en == 1) begin
				if(push == 1) begin
					count	<=	count + 1;
				end
			end
			else begin
				count	<=	2'd3;
			end
		end
	end

	always @(`CLK_RST_EDGE)
		if (`RST)			cnt_en <= 0;
		else if (push)			cnt_en <= 1;
		else if (end_cnt_en)		cnt_en <= 0;

	always @(`CLK_RST_EDGE)
		if (`RST)	cnt <= 0;
		else if(cnt_en)	cnt <= cnt_max? 0: cnt + 1;

	always @(`CLK_RST_EDGE)
		if (`RST)	ready <= 0;
		else 		ready <= cnt_en;

	always @(posedge clk) begin
		if (cnt_en == 1'b0) begin
			dt	<=	1'b0;
		end
		else	begin	//1) W_1(66), 2) D_3(167), 3) N_13(166), 4) P_15(1666)
			case	(count)
				2'd0	:	begin
					case (cnt)
						10'd0	:	dt	<=	92	;
						10'd1	:	dt	<=	101	;
						10'd2	:	dt	<=	84	;
						10'd3	:	dt	<=	67	;
						10'd4	:	dt	<=	68	;
						10'd5	:	dt	<=	58	;
						10'd6	:	dt	<=	73	;
						10'd7	:	dt	<=	20	;
						10'd8	:	dt	<=	55	;
						10'd9	:	dt	<=	85	;
						10'd10	:	dt	<=	98	;
						10'd11	:	dt	<=	108	;
						10'd12	:	dt	<=	150	;
						10'd13	:	dt	<=	117	;
						10'd14	:	dt	<=	99	;
						10'd15	:	dt	<=	136	;
						10'd16	:	dt	<=	135	;
						10'd17	:	dt	<=	142	;
						10'd18	:	dt	<=	143	;
						10'd19	:	dt	<=	146	;
						10'd20	:	dt	<=	150	;
						10'd21	:	dt	<=	153	;
						10'd22	:	dt	<=	154	;
						10'd23	:	dt	<=	157	;
						10'd24	:	dt	<=	158	;
						10'd25	:	dt	<=	160	;
						10'd26	:	dt	<=	162	;
						10'd27	:	dt	<=	163	;
						10'd28	:	dt	<=	95	;
						10'd29	:	dt	<=	104	;
						10'd30	:	dt	<=	82	;
						10'd31	:	dt	<=	71	;
						10'd32	:	dt	<=	66	;
						10'd33	:	dt	<=	65	;
						10'd34	:	dt	<=	71	;
						10'd35	:	dt	<=	20	;
						10'd36	:	dt	<=	62	;
						10'd37	:	dt	<=	87	;
						10'd38	:	dt	<=	104	;
						10'd39	:	dt	<=	112	;
						10'd40	:	dt	<=	152	;
						10'd41	:	dt	<=	130	;
						10'd42	:	dt	<=	85	;
						10'd43	:	dt	<=	136	;
						10'd44	:	dt	<=	105	;
						10'd45	:	dt	<=	132	;
						10'd46	:	dt	<=	148	;
						10'd47	:	dt	<=	148	;
						10'd48	:	dt	<=	151	;
						10'd49	:	dt	<=	154	;
						10'd50	:	dt	<=	156	;
						10'd51	:	dt	<=	160	;
						10'd52	:	dt	<=	160	;
						10'd53	:	dt	<=	162	;
						10'd54	:	dt	<=	163	;
						10'd55	:	dt	<=	164	;
						10'd56	:	dt	<=	97	;
						10'd57	:	dt	<=	106	;
						10'd58	:	dt	<=	79	;
						10'd59	:	dt	<=	74	;
						10'd60	:	dt	<=	63	;
						10'd61	:	dt	<=	72	;
						10'd62	:	dt	<=	65	;
						10'd63	:	dt	<=	22	;
						10'd64	:	dt	<=	69	;
						10'd65	:	dt	<=	84	;
						10'd66	:	dt	<=	140	;
						10'd67	:	dt	<=	122	;
						10'd68	:	dt	<=	123	;
						10'd69	:	dt	<=	151	;
						10'd70	:	dt	<=	95	;
						10'd71	:	dt	<=	148	;
						10'd72	:	dt	<=	103	;
						10'd73	:	dt	<=	101	;
						10'd74	:	dt	<=	153	;
						10'd75	:	dt	<=	148	;
						10'd76	:	dt	<=	153	;
						10'd77	:	dt	<=	154	;
						10'd78	:	dt	<=	158	;
						10'd79	:	dt	<=	160	;
						10'd80	:	dt	<=	161	;
						10'd81	:	dt	<=	162	;
						10'd82	:	dt	<=	163	;
						10'd83	:	dt	<=	165	;
						10'd84	:	dt	<=	101	;
						10'd85	:	dt	<=	106	;
						10'd86	:	dt	<=	76	;
						10'd87	:	dt	<=	78	;
						10'd88	:	dt	<=	64	;
						10'd89	:	dt	<=	79	;
						10'd90	:	dt	<=	56	;
						10'd91	:	dt	<=	25	;
						10'd92	:	dt	<=	73	;
						10'd93	:	dt	<=	86	;
						10'd94	:	dt	<=	151	;
						10'd95	:	dt	<=	131	;
						10'd96	:	dt	<=	110	;
						10'd97	:	dt	<=	154	;
						10'd98	:	dt	<=	100	;
						10'd99	:	dt	<=	150	;
						10'd100	:	dt	<=	131	;
						10'd101	:	dt	<=	88	;
						10'd102	:	dt	<=	149	;
						10'd103	:	dt	<=	152	;
						10'd104	:	dt	<=	154	;
						10'd105	:	dt	<=	156	;
						10'd106	:	dt	<=	159	;
						10'd107	:	dt	<=	161	;
						10'd108	:	dt	<=	162	;
						10'd109	:	dt	<=	164	;
						10'd110	:	dt	<=	165	;
						10'd111	:	dt	<=	166	;
						10'd112	:	dt	<=	104	;
						10'd113	:	dt	<=	104	;
						10'd114	:	dt	<=	75	;
						10'd115	:	dt	<=	81	;
						10'd116	:	dt	<=	62	;
						10'd117	:	dt	<=	84	;
						10'd118	:	dt	<=	47	;
						10'd119	:	dt	<=	31	;
						10'd120	:	dt	<=	79	;
						10'd121	:	dt	<=	89	;
						10'd122	:	dt	<=	153	;
						10'd123	:	dt	<=	138	;
						10'd124	:	dt	<=	110	;
						10'd125	:	dt	<=	170	;
						10'd126	:	dt	<=	124	;
						10'd127	:	dt	<=	135	;
						10'd128	:	dt	<=	144	;
						10'd129	:	dt	<=	87	;
						10'd130	:	dt	<=	140	;
						10'd131	:	dt	<=	156	;
						10'd132	:	dt	<=	154	;
						10'd133	:	dt	<=	158	;
						10'd134	:	dt	<=	160	;
						10'd135	:	dt	<=	162	;
						10'd136	:	dt	<=	164	;
						10'd137	:	dt	<=	166	;
						10'd138	:	dt	<=	168	;
						10'd139	:	dt	<=	168	;
						10'd140	:	dt	<=	108	;
						10'd141	:	dt	<=	103	;
						10'd142	:	dt	<=	78	;
						10'd143	:	dt	<=	84	;
						10'd144	:	dt	<=	64	;
						10'd145	:	dt	<=	89	;
						10'd146	:	dt	<=	38	;
						10'd147	:	dt	<=	39	;
						10'd148	:	dt	<=	81	;
						10'd149	:	dt	<=	89	;
						10'd150	:	dt	<=	152	;
						10'd151	:	dt	<=	144	;
						10'd152	:	dt	<=	111	;
						10'd153	:	dt	<=	179	;
						10'd154	:	dt	<=	133	;
						10'd155	:	dt	<=	129	;
						10'd156	:	dt	<=	166	;
						10'd157	:	dt	<=	100	;
						10'd158	:	dt	<=	126	;
						10'd159	:	dt	<=	161	;
						10'd160	:	dt	<=	157	;
						10'd161	:	dt	<=	160	;
						10'd162	:	dt	<=	162	;
						10'd163	:	dt	<=	164	;
						10'd164	:	dt	<=	166	;
						10'd165	:	dt	<=	169	;
						10'd166	:	dt	<=	170	;
						10'd167	:	dt	<=	170	;
						10'd168	:	dt	<=	112	;
						10'd169	:	dt	<=	100	;
						10'd170	:	dt	<=	82	;
						10'd171	:	dt	<=	88	;
						10'd172	:	dt	<=	66	;
						10'd173	:	dt	<=	93	;
						10'd174	:	dt	<=	32	;
						10'd175	:	dt	<=	42	;
						10'd176	:	dt	<=	111	;
						10'd177	:	dt	<=	112	;
						10'd178	:	dt	<=	145	;
						10'd179	:	dt	<=	166	;
						10'd180	:	dt	<=	116	;
						10'd181	:	dt	<=	169	;
						10'd182	:	dt	<=	136	;
						10'd183	:	dt	<=	133	;
						10'd184	:	dt	<=	179	;
						10'd185	:	dt	<=	117	;
						10'd186	:	dt	<=	108	;
						10'd187	:	dt	<=	163	;
						10'd188	:	dt	<=	159	;
						10'd189	:	dt	<=	162	;
						10'd190	:	dt	<=	164	;
						10'd191	:	dt	<=	167	;
						10'd192	:	dt	<=	170	;
						10'd193	:	dt	<=	171	;
						10'd194	:	dt	<=	171	;
						10'd195	:	dt	<=	172	;
						10'd196	:	dt	<=	115	;
						10'd197	:	dt	<=	99	;
						10'd198	:	dt	<=	86	;
						10'd199	:	dt	<=	86	;
						10'd200	:	dt	<=	69	;
						10'd201	:	dt	<=	94	;
						10'd202	:	dt	<=	27	;
						10'd203	:	dt	<=	49	;
						10'd204	:	dt	<=	149	;
						10'd205	:	dt	<=	119	;
						10'd206	:	dt	<=	136	;
						10'd207	:	dt	<=	169	;
						10'd208	:	dt	<=	114	;
						10'd209	:	dt	<=	158	;
						10'd210	:	dt	<=	141	;
						10'd211	:	dt	<=	124	;
						10'd212	:	dt	<=	173	;
						10'd213	:	dt	<=	130	;
						10'd214	:	dt	<=	100	;
						10'd215	:	dt	<=	161	;
						10'd216	:	dt	<=	161	;
						10'd217	:	dt	<=	162	;
						10'd218	:	dt	<=	166	;
						10'd219	:	dt	<=	169	;
						10'd220	:	dt	<=	171	;
						10'd221	:	dt	<=	172	;
						10'd222	:	dt	<=	172	;
						10'd223	:	dt	<=	173	;
						10'd224	:	dt	<=	118	;
						10'd225	:	dt	<=	97	;
						10'd226	:	dt	<=	89	;
						10'd227	:	dt	<=	84	;
						10'd228	:	dt	<=	75	;
						10'd229	:	dt	<=	91	;
						10'd230	:	dt	<=	23	;
						10'd231	:	dt	<=	59	;
						10'd232	:	dt	<=	152	;
						10'd233	:	dt	<=	114	;
						10'd234	:	dt	<=	132	;
						10'd235	:	dt	<=	168	;
						10'd236	:	dt	<=	110	;
						10'd237	:	dt	<=	156	;
						10'd238	:	dt	<=	156	;
						10'd239	:	dt	<=	117	;
						10'd240	:	dt	<=	169	;
						10'd241	:	dt	<=	139	;
						10'd242	:	dt	<=	98	;
						10'd243	:	dt	<=	160	;
						10'd244	:	dt	<=	163	;
						10'd245	:	dt	<=	165	;
						10'd246	:	dt	<=	169	;
						10'd247	:	dt	<=	171	;
						10'd248	:	dt	<=	172	;
						10'd249	:	dt	<=	174	;
						10'd250	:	dt	<=	175	;
						10'd251	:	dt	<=	176	;
						10'd252	:	dt	<=	118	;
						10'd253	:	dt	<=	95	;
						10'd254	:	dt	<=	93	;
						10'd255	:	dt	<=	82	;
						10'd256	:	dt	<=	81	;
						10'd257	:	dt	<=	87	;
						10'd258	:	dt	<=	22	;
						10'd259	:	dt	<=	64	;
						10'd260	:	dt	<=	157	;
						10'd261	:	dt	<=	118	;
						10'd262	:	dt	<=	126	;
						10'd263	:	dt	<=	176	;
						10'd264	:	dt	<=	110	;
						10'd265	:	dt	<=	150	;
						10'd266	:	dt	<=	168	;
						10'd267	:	dt	<=	114	;
						10'd268	:	dt	<=	174	;
						10'd269	:	dt	<=	149	;
						10'd270	:	dt	<=	99	;
						10'd271	:	dt	<=	155	;
						10'd272	:	dt	<=	165	;
						10'd273	:	dt	<=	168	;
						10'd274	:	dt	<=	170	;
						10'd275	:	dt	<=	173	;
						10'd276	:	dt	<=	174	;
						10'd277	:	dt	<=	176	;
						10'd278	:	dt	<=	177	;
						10'd279	:	dt	<=	176	;
						10'd280	:	dt	<=	119	;
						10'd281	:	dt	<=	94	;
						10'd282	:	dt	<=	98	;
						10'd283	:	dt	<=	80	;
						10'd284	:	dt	<=	89	;
						10'd285	:	dt	<=	78	;
						10'd286	:	dt	<=	24	;
						10'd287	:	dt	<=	67	;
						10'd288	:	dt	<=	163	;
						10'd289	:	dt	<=	139	;
						10'd290	:	dt	<=	123	;
						10'd291	:	dt	<=	180	;
						10'd292	:	dt	<=	120	;
						10'd293	:	dt	<=	127	;
						10'd294	:	dt	<=	170	;
						10'd295	:	dt	<=	107	;
						10'd296	:	dt	<=	161	;
						10'd297	:	dt	<=	153	;
						10'd298	:	dt	<=	94	;
						10'd299	:	dt	<=	148	;
						10'd300	:	dt	<=	171	;
						10'd301	:	dt	<=	169	;
						10'd302	:	dt	<=	171	;
						10'd303	:	dt	<=	174	;
						10'd304	:	dt	<=	176	;
						10'd305	:	dt	<=	177	;
						10'd306	:	dt	<=	177	;
						10'd307	:	dt	<=	177	;
						10'd308	:	dt	<=	115	;
						10'd309	:	dt	<=	95	;
						10'd310	:	dt	<=	102	;
						10'd311	:	dt	<=	78	;
						10'd312	:	dt	<=	97	;
						10'd313	:	dt	<=	68	;
						10'd314	:	dt	<=	28	;
						10'd315	:	dt	<=	70	;
						10'd316	:	dt	<=	158	;
						10'd317	:	dt	<=	142	;
						10'd318	:	dt	<=	107	;
						10'd319	:	dt	<=	179	;
						10'd320	:	dt	<=	126	;
						10'd321	:	dt	<=	98	;
						10'd322	:	dt	<=	161	;
						10'd323	:	dt	<=	99	;
						10'd324	:	dt	<=	143	;
						10'd325	:	dt	<=	163	;
						10'd326	:	dt	<=	95	;
						10'd327	:	dt	<=	140	;
						10'd328	:	dt	<=	174	;
						10'd329	:	dt	<=	168	;
						10'd330	:	dt	<=	172	;
						10'd331	:	dt	<=	176	;
						10'd332	:	dt	<=	177	;
						10'd333	:	dt	<=	178	;
						10'd334	:	dt	<=	179	;
						10'd335	:	dt	<=	178	;
						10'd336	:	dt	<=	114	;
						10'd337	:	dt	<=	96	;
						10'd338	:	dt	<=	103	;
						10'd339	:	dt	<=	75	;
						10'd340	:	dt	<=	103	;
						10'd341	:	dt	<=	58	;
						10'd342	:	dt	<=	33	;
						10'd343	:	dt	<=	72	;
						10'd344	:	dt	<=	146	;
						10'd345	:	dt	<=	149	;
						10'd346	:	dt	<=	100	;
						10'd347	:	dt	<=	161	;
						10'd348	:	dt	<=	136	;
						10'd349	:	dt	<=	128	;
						10'd350	:	dt	<=	148	;
						10'd351	:	dt	<=	141	;
						10'd352	:	dt	<=	157	;
						10'd353	:	dt	<=	139	;
						10'd354	:	dt	<=	91	;
						10'd355	:	dt	<=	122	;
						10'd356	:	dt	<=	176	;
						10'd357	:	dt	<=	169	;
						10'd358	:	dt	<=	174	;
						10'd359	:	dt	<=	176	;
						10'd360	:	dt	<=	178	;
						10'd361	:	dt	<=	180	;
						10'd362	:	dt	<=	180	;
						10'd363	:	dt	<=	179	;
						10'd364	:	dt	<=	113	;
						10'd365	:	dt	<=	96	;
						10'd366	:	dt	<=	103	;
						10'd367	:	dt	<=	74	;
						10'd368	:	dt	<=	108	;
						10'd369	:	dt	<=	48	;
						10'd370	:	dt	<=	39	;
						10'd371	:	dt	<=	74	;
						10'd372	:	dt	<=	143	;
						10'd373	:	dt	<=	166	;
						10'd374	:	dt	<=	100	;
						10'd375	:	dt	<=	142	;
						10'd376	:	dt	<=	160	;
						10'd377	:	dt	<=	137	;
						10'd378	:	dt	<=	121	;
						10'd379	:	dt	<=	154	;
						10'd380	:	dt	<=	155	;
						10'd381	:	dt	<=	103	;
						10'd382	:	dt	<=	78	;
						10'd383	:	dt	<=	107	;
						10'd384	:	dt	<=	177	;
						10'd385	:	dt	<=	172	;
						10'd386	:	dt	<=	175	;
						10'd387	:	dt	<=	177	;
						10'd388	:	dt	<=	179	;
						10'd389	:	dt	<=	180	;
						10'd390	:	dt	<=	181	;
						10'd391	:	dt	<=	183	;
						10'd392	:	dt	<=	110	;
						10'd393	:	dt	<=	99	;
						10'd394	:	dt	<=	103	;
						10'd395	:	dt	<=	73	;
						10'd396	:	dt	<=	111	;
						10'd397	:	dt	<=	39	;
						10'd398	:	dt	<=	45	;
						10'd399	:	dt	<=	76	;
						10'd400	:	dt	<=	144	;
						10'd401	:	dt	<=	155	;
						10'd402	:	dt	<=	122	;
						10'd403	:	dt	<=	152	;
						10'd404	:	dt	<=	152	;
						10'd405	:	dt	<=	150	;
						10'd406	:	dt	<=	142	;
						10'd407	:	dt	<=	178	;
						10'd408	:	dt	<=	168	;
						10'd409	:	dt	<=	110	;
						10'd410	:	dt	<=	72	;
						10'd411	:	dt	<=	87	;
						10'd412	:	dt	<=	170	;
						10'd413	:	dt	<=	174	;
						10'd414	:	dt	<=	177	;
						10'd415	:	dt	<=	179	;
						10'd416	:	dt	<=	180	;
						10'd417	:	dt	<=	181	;
						10'd418	:	dt	<=	183	;
						10'd419	:	dt	<=	184	;
						10'd420	:	dt	<=	109	;
						10'd421	:	dt	<=	103	;
						10'd422	:	dt	<=	102	;
						10'd423	:	dt	<=	74	;
						10'd424	:	dt	<=	111	;
						10'd425	:	dt	<=	31	;
						10'd426	:	dt	<=	51	;
						10'd427	:	dt	<=	78	;
						10'd428	:	dt	<=	146	;
						10'd429	:	dt	<=	160	;
						10'd430	:	dt	<=	159	;
						10'd431	:	dt	<=	142	;
						10'd432	:	dt	<=	141	;
						10'd433	:	dt	<=	146	;
						10'd434	:	dt	<=	154	;
						10'd435	:	dt	<=	168	;
						10'd436	:	dt	<=	161	;
						10'd437	:	dt	<=	136	;
						10'd438	:	dt	<=	89	;
						10'd439	:	dt	<=	67	;
						10'd440	:	dt	<=	159	;
						10'd441	:	dt	<=	178	;
						10'd442	:	dt	<=	176	;
						10'd443	:	dt	<=	179	;
						10'd444	:	dt	<=	180	;
						10'd445	:	dt	<=	182	;
						10'd446	:	dt	<=	182	;
						10'd447	:	dt	<=	184	;
						10'd448	:	dt	<=	108	;
						10'd449	:	dt	<=	105	;
						10'd450	:	dt	<=	100	;
						10'd451	:	dt	<=	80	;
						10'd452	:	dt	<=	111	;
						10'd453	:	dt	<=	24	;
						10'd454	:	dt	<=	57	;
						10'd455	:	dt	<=	79	;
						10'd456	:	dt	<=	160	;
						10'd457	:	dt	<=	178	;
						10'd458	:	dt	<=	151	;
						10'd459	:	dt	<=	129	;
						10'd460	:	dt	<=	128	;
						10'd461	:	dt	<=	133	;
						10'd462	:	dt	<=	139	;
						10'd463	:	dt	<=	136	;
						10'd464	:	dt	<=	158	;
						10'd465	:	dt	<=	162	;
						10'd466	:	dt	<=	122	;
						10'd467	:	dt	<=	69	;
						10'd468	:	dt	<=	141	;
						10'd469	:	dt	<=	183	;
						10'd470	:	dt	<=	176	;
						10'd471	:	dt	<=	180	;
						10'd472	:	dt	<=	180	;
						10'd473	:	dt	<=	182	;
						10'd474	:	dt	<=	183	;
						10'd475	:	dt	<=	185	;
						10'd476	:	dt	<=	105	;
						10'd477	:	dt	<=	111	;
						10'd478	:	dt	<=	97	;
						10'd479	:	dt	<=	87	;
						10'd480	:	dt	<=	107	;
						10'd481	:	dt	<=	20	;
						10'd482	:	dt	<=	60	;
						10'd483	:	dt	<=	82	;
						10'd484	:	dt	<=	168	;
						10'd485	:	dt	<=	172	;
						10'd486	:	dt	<=	138	;
						10'd487	:	dt	<=	119	;
						10'd488	:	dt	<=	127	;
						10'd489	:	dt	<=	137	;
						10'd490	:	dt	<=	152	;
						10'd491	:	dt	<=	167	;
						10'd492	:	dt	<=	171	;
						10'd493	:	dt	<=	178	;
						10'd494	:	dt	<=	154	;
						10'd495	:	dt	<=	91	;
						10'd496	:	dt	<=	114	;
						10'd497	:	dt	<=	183	;
						10'd498	:	dt	<=	177	;
						10'd499	:	dt	<=	180	;
						10'd500	:	dt	<=	181	;
						10'd501	:	dt	<=	183	;
						10'd502	:	dt	<=	184	;
						10'd503	:	dt	<=	184	;
						10'd504	:	dt	<=	104	;
						10'd505	:	dt	<=	114	;
						10'd506	:	dt	<=	94	;
						10'd507	:	dt	<=	94	;
						10'd508	:	dt	<=	101	;
						10'd509	:	dt	<=	19	;
						10'd510	:	dt	<=	65	;
						10'd511	:	dt	<=	82	;
						10'd512	:	dt	<=	156	;
						10'd513	:	dt	<=	171	;
						10'd514	:	dt	<=	131	;
						10'd515	:	dt	<=	115	;
						10'd516	:	dt	<=	135	;
						10'd517	:	dt	<=	137	;
						10'd518	:	dt	<=	160	;
						10'd519	:	dt	<=	191	;
						10'd520	:	dt	<=	176	;
						10'd521	:	dt	<=	179	;
						10'd522	:	dt	<=	165	;
						10'd523	:	dt	<=	114	;
						10'd524	:	dt	<=	96	;
						10'd525	:	dt	<=	180	;
						10'd526	:	dt	<=	177	;
						10'd527	:	dt	<=	180	;
						10'd528	:	dt	<=	181	;
						10'd529	:	dt	<=	183	;
						10'd530	:	dt	<=	184	;
						10'd531	:	dt	<=	184	;
						10'd532	:	dt	<=	107	;
						10'd533	:	dt	<=	116	;
						10'd534	:	dt	<=	90	;
						10'd535	:	dt	<=	100	;
						10'd536	:	dt	<=	91	;
						10'd537	:	dt	<=	19	;
						10'd538	:	dt	<=	71	;
						10'd539	:	dt	<=	82	;
						10'd540	:	dt	<=	137	;
						10'd541	:	dt	<=	176	;
						10'd542	:	dt	<=	141	;
						10'd543	:	dt	<=	122	;
						10'd544	:	dt	<=	128	;
						10'd545	:	dt	<=	145	;
						10'd546	:	dt	<=	164	;
						10'd547	:	dt	<=	190	;
						10'd548	:	dt	<=	186	;
						10'd549	:	dt	<=	169	;
						10'd550	:	dt	<=	153	;
						10'd551	:	dt	<=	110	;
						10'd552	:	dt	<=	94	;
						10'd553	:	dt	<=	179	;
						10'd554	:	dt	<=	178	;
						10'd555	:	dt	<=	181	;
						10'd556	:	dt	<=	182	;
						10'd557	:	dt	<=	184	;
						10'd558	:	dt	<=	185	;
						10'd559	:	dt	<=	186	;
						10'd560	:	dt	<=	107	;
						10'd561	:	dt	<=	117	;
						10'd562	:	dt	<=	86	;
						10'd563	:	dt	<=	107	;
						10'd564	:	dt	<=	82	;
						10'd565	:	dt	<=	20	;
						10'd566	:	dt	<=	73	;
						10'd567	:	dt	<=	85	;
						10'd568	:	dt	<=	115	;
						10'd569	:	dt	<=	173	;
						10'd570	:	dt	<=	148	;
						10'd571	:	dt	<=	129	;
						10'd572	:	dt	<=	125	;
						10'd573	:	dt	<=	151	;
						10'd574	:	dt	<=	166	;
						10'd575	:	dt	<=	192	;
						10'd576	:	dt	<=	188	;
						10'd577	:	dt	<=	166	;
						10'd578	:	dt	<=	142	;
						10'd579	:	dt	<=	96	;
						10'd580	:	dt	<=	101	;
						10'd581	:	dt	<=	183	;
						10'd582	:	dt	<=	177	;
						10'd583	:	dt	<=	180	;
						10'd584	:	dt	<=	183	;
						10'd585	:	dt	<=	184	;
						10'd586	:	dt	<=	185	;
						10'd587	:	dt	<=	186	;
						10'd588	:	dt	<=	107	;
						10'd589	:	dt	<=	119	;
						10'd590	:	dt	<=	84	;
						10'd591	:	dt	<=	114	;
						10'd592	:	dt	<=	73	;
						10'd593	:	dt	<=	22	;
						10'd594	:	dt	<=	74	;
						10'd595	:	dt	<=	89	;
						10'd596	:	dt	<=	101	;
						10'd597	:	dt	<=	160	;
						10'd598	:	dt	<=	163	;
						10'd599	:	dt	<=	138	;
						10'd600	:	dt	<=	123	;
						10'd601	:	dt	<=	144	;
						10'd602	:	dt	<=	164	;
						10'd603	:	dt	<=	188	;
						10'd604	:	dt	<=	184	;
						10'd605	:	dt	<=	161	;
						10'd606	:	dt	<=	138	;
						10'd607	:	dt	<=	92	;
						10'd608	:	dt	<=	104	;
						10'd609	:	dt	<=	184	;
						10'd610	:	dt	<=	177	;
						10'd611	:	dt	<=	180	;
						10'd612	:	dt	<=	183	;
						10'd613	:	dt	<=	185	;
						10'd614	:	dt	<=	185	;
						10'd615	:	dt	<=	186	;
						10'd616	:	dt	<=	111	;
						10'd617	:	dt	<=	122	;
						10'd618	:	dt	<=	82	;
						10'd619	:	dt	<=	123	;
						10'd620	:	dt	<=	64	;
						10'd621	:	dt	<=	26	;
						10'd622	:	dt	<=	75	;
						10'd623	:	dt	<=	89	;
						10'd624	:	dt	<=	96	;
						10'd625	:	dt	<=	144	;
						10'd626	:	dt	<=	170	;
						10'd627	:	dt	<=	147	;
						10'd628	:	dt	<=	134	;
						10'd629	:	dt	<=	133	;
						10'd630	:	dt	<=	158	;
						10'd631	:	dt	<=	183	;
						10'd632	:	dt	<=	175	;
						10'd633	:	dt	<=	153	;
						10'd634	:	dt	<=	136	;
						10'd635	:	dt	<=	89	;
						10'd636	:	dt	<=	104	;
						10'd637	:	dt	<=	183	;
						10'd638	:	dt	<=	178	;
						10'd639	:	dt	<=	182	;
						10'd640	:	dt	<=	184	;
						10'd641	:	dt	<=	184	;
						10'd642	:	dt	<=	185	;
						10'd643	:	dt	<=	186	;
						10'd644	:	dt	<=	115	;
						10'd645	:	dt	<=	124	;
						10'd646	:	dt	<=	81	;
						10'd647	:	dt	<=	131	;
						10'd648	:	dt	<=	55	;
						10'd649	:	dt	<=	30	;
						10'd650	:	dt	<=	77	;
						10'd651	:	dt	<=	88	;
						10'd652	:	dt	<=	98	;
						10'd653	:	dt	<=	119	;
						10'd654	:	dt	<=	162	;
						10'd655	:	dt	<=	155	;
						10'd656	:	dt	<=	148	;
						10'd657	:	dt	<=	134	;
						10'd658	:	dt	<=	150	;
						10'd659	:	dt	<=	176	;
						10'd660	:	dt	<=	166	;
						10'd661	:	dt	<=	145	;
						10'd662	:	dt	<=	129	;
						10'd663	:	dt	<=	85	;
						10'd664	:	dt	<=	110	;
						10'd665	:	dt	<=	184	;
						10'd666	:	dt	<=	178	;
						10'd667	:	dt	<=	183	;
						10'd668	:	dt	<=	184	;
						10'd669	:	dt	<=	184	;
						10'd670	:	dt	<=	185	;
						10'd671	:	dt	<=	185	;
						10'd672	:	dt	<=	120	;
						10'd673	:	dt	<=	124	;
						10'd674	:	dt	<=	84	;
						10'd675	:	dt	<=	134	;
						10'd676	:	dt	<=	45	;
						10'd677	:	dt	<=	34	;
						10'd678	:	dt	<=	75	;
						10'd679	:	dt	<=	86	;
						10'd680	:	dt	<=	98	;
						10'd681	:	dt	<=	107	;
						10'd682	:	dt	<=	139	;
						10'd683	:	dt	<=	161	;
						10'd684	:	dt	<=	153	;
						10'd685	:	dt	<=	145	;
						10'd686	:	dt	<=	140	;
						10'd687	:	dt	<=	157	;
						10'd688	:	dt	<=	160	;
						10'd689	:	dt	<=	138	;
						10'd690	:	dt	<=	124	;
						10'd691	:	dt	<=	82	;
						10'd692	:	dt	<=	126	;
						10'd693	:	dt	<=	182	;
						10'd694	:	dt	<=	176	;
						10'd695	:	dt	<=	180	;
						10'd696	:	dt	<=	181	;
						10'd697	:	dt	<=	182	;
						10'd698	:	dt	<=	183	;
						10'd699	:	dt	<=	183	;
						10'd700	:	dt	<=	124	;
						10'd701	:	dt	<=	121	;
						10'd702	:	dt	<=	86	;
						10'd703	:	dt	<=	136	;
						10'd704	:	dt	<=	36	;
						10'd705	:	dt	<=	38	;
						10'd706	:	dt	<=	72	;
						10'd707	:	dt	<=	84	;
						10'd708	:	dt	<=	95	;
						10'd709	:	dt	<=	106	;
						10'd710	:	dt	<=	118	;
						10'd711	:	dt	<=	156	;
						10'd712	:	dt	<=	156	;
						10'd713	:	dt	<=	148	;
						10'd714	:	dt	<=	132	;
						10'd715	:	dt	<=	135	;
						10'd716	:	dt	<=	148	;
						10'd717	:	dt	<=	126	;
						10'd718	:	dt	<=	115	;
						10'd719	:	dt	<=	85	;
						10'd720	:	dt	<=	150	;
						10'd721	:	dt	<=	179	;
						10'd722	:	dt	<=	175	;
						10'd723	:	dt	<=	178	;
						10'd724	:	dt	<=	179	;
						10'd725	:	dt	<=	180	;
						10'd726	:	dt	<=	182	;
						10'd727	:	dt	<=	182	;
						10'd728	:	dt	<=	126	;
						10'd729	:	dt	<=	116	;
						10'd730	:	dt	<=	90	;
						10'd731	:	dt	<=	136	;
						10'd732	:	dt	<=	27	;
						10'd733	:	dt	<=	41	;
						10'd734	:	dt	<=	71	;
						10'd735	:	dt	<=	81	;
						10'd736	:	dt	<=	93	;
						10'd737	:	dt	<=	107	;
						10'd738	:	dt	<=	109	;
						10'd739	:	dt	<=	148	;
						10'd740	:	dt	<=	157	;
						10'd741	:	dt	<=	141	;
						10'd742	:	dt	<=	127	;
						10'd743	:	dt	<=	126	;
						10'd744	:	dt	<=	127	;
						10'd745	:	dt	<=	121	;
						10'd746	:	dt	<=	113	;
						10'd747	:	dt	<=	85	;
						10'd748	:	dt	<=	161	;
						10'd749	:	dt	<=	173	;
						10'd750	:	dt	<=	173	;
						10'd751	:	dt	<=	177	;
						10'd752	:	dt	<=	179	;
						10'd753	:	dt	<=	180	;
						10'd754	:	dt	<=	182	;
						10'd755	:	dt	<=	182	;
						10'd756	:	dt	<=	130	;
						10'd757	:	dt	<=	113	;
						10'd758	:	dt	<=	94	;
						10'd759	:	dt	<=	130	;
						10'd760	:	dt	<=	25	;
						10'd761	:	dt	<=	45	;
						10'd762	:	dt	<=	68	;
						10'd763	:	dt	<=	74	;
						10'd764	:	dt	<=	85	;
						10'd765	:	dt	<=	100	;
						10'd766	:	dt	<=	103	;
						10'd767	:	dt	<=	139	;
						10'd768	:	dt	<=	152	;
						10'd769	:	dt	<=	130	;
						10'd770	:	dt	<=	129	;
						10'd771	:	dt	<=	134	;
						10'd772	:	dt	<=	128	;
						10'd773	:	dt	<=	121	;
						10'd774	:	dt	<=	106	;
						10'd775	:	dt	<=	81	;
						10'd776	:	dt	<=	162	;
						10'd777	:	dt	<=	170	;
						10'd778	:	dt	<=	170	;
						10'd779	:	dt	<=	174	;
						10'd780	:	dt	<=	176	;
						10'd781	:	dt	<=	178	;
						10'd782	:	dt	<=	179	;
						10'd783	:	dt	<=	178	;

					endcase
				end
				2'd1	:	begin
					case (cnt)
						10'd0	:	dt	<=	132	;
						10'd1	:	dt	<=	135	;
						10'd2	:	dt	<=	135	;
						10'd3	:	dt	<=	135	;
						10'd4	:	dt	<=	135	;
						10'd5	:	dt	<=	136	;
						10'd6	:	dt	<=	137	;
						10'd7	:	dt	<=	136	;
						10'd8	:	dt	<=	137	;
						10'd9	:	dt	<=	136	;
						10'd10	:	dt	<=	136	;
						10'd11	:	dt	<=	136	;
						10'd12	:	dt	<=	135	;
						10'd13	:	dt	<=	134	;
						10'd14	:	dt	<=	132	;
						10'd15	:	dt	<=	131	;
						10'd16	:	dt	<=	129	;
						10'd17	:	dt	<=	121	;
						10'd18	:	dt	<=	130	;
						10'd19	:	dt	<=	126	;
						10'd20	:	dt	<=	126	;
						10'd21	:	dt	<=	125	;
						10'd22	:	dt	<=	122	;
						10'd23	:	dt	<=	121	;
						10'd24	:	dt	<=	118	;
						10'd25	:	dt	<=	117	;
						10'd26	:	dt	<=	115	;
						10'd27	:	dt	<=	113	;
						10'd28	:	dt	<=	136	;
						10'd29	:	dt	<=	138	;
						10'd30	:	dt	<=	138	;
						10'd31	:	dt	<=	139	;
						10'd32	:	dt	<=	138	;
						10'd33	:	dt	<=	138	;
						10'd34	:	dt	<=	139	;
						10'd35	:	dt	<=	140	;
						10'd36	:	dt	<=	139	;
						10'd37	:	dt	<=	139	;
						10'd38	:	dt	<=	141	;
						10'd39	:	dt	<=	140	;
						10'd40	:	dt	<=	138	;
						10'd41	:	dt	<=	137	;
						10'd42	:	dt	<=	136	;
						10'd43	:	dt	<=	135	;
						10'd44	:	dt	<=	141	;
						10'd45	:	dt	<=	77	;
						10'd46	:	dt	<=	108	;
						10'd47	:	dt	<=	136	;
						10'd48	:	dt	<=	129	;
						10'd49	:	dt	<=	127	;
						10'd50	:	dt	<=	126	;
						10'd51	:	dt	<=	125	;
						10'd52	:	dt	<=	122	;
						10'd53	:	dt	<=	121	;
						10'd54	:	dt	<=	118	;
						10'd55	:	dt	<=	116	;
						10'd56	:	dt	<=	139	;
						10'd57	:	dt	<=	142	;
						10'd58	:	dt	<=	142	;
						10'd59	:	dt	<=	142	;
						10'd60	:	dt	<=	143	;
						10'd61	:	dt	<=	143	;
						10'd62	:	dt	<=	143	;
						10'd63	:	dt	<=	144	;
						10'd64	:	dt	<=	143	;
						10'd65	:	dt	<=	143	;
						10'd66	:	dt	<=	144	;
						10'd67	:	dt	<=	145	;
						10'd68	:	dt	<=	143	;
						10'd69	:	dt	<=	142	;
						10'd70	:	dt	<=	140	;
						10'd71	:	dt	<=	140	;
						10'd72	:	dt	<=	132	;
						10'd73	:	dt	<=	58	;
						10'd74	:	dt	<=	77	;
						10'd75	:	dt	<=	145	;
						10'd76	:	dt	<=	131	;
						10'd77	:	dt	<=	131	;
						10'd78	:	dt	<=	130	;
						10'd79	:	dt	<=	129	;
						10'd80	:	dt	<=	127	;
						10'd81	:	dt	<=	124	;
						10'd82	:	dt	<=	122	;
						10'd83	:	dt	<=	119	;
						10'd84	:	dt	<=	144	;
						10'd85	:	dt	<=	145	;
						10'd86	:	dt	<=	146	;
						10'd87	:	dt	<=	145	;
						10'd88	:	dt	<=	147	;
						10'd89	:	dt	<=	147	;
						10'd90	:	dt	<=	148	;
						10'd91	:	dt	<=	149	;
						10'd92	:	dt	<=	149	;
						10'd93	:	dt	<=	148	;
						10'd94	:	dt	<=	147	;
						10'd95	:	dt	<=	146	;
						10'd96	:	dt	<=	147	;
						10'd97	:	dt	<=	146	;
						10'd98	:	dt	<=	144	;
						10'd99	:	dt	<=	143	;
						10'd100	:	dt	<=	131	;
						10'd101	:	dt	<=	56	;
						10'd102	:	dt	<=	58	;
						10'd103	:	dt	<=	146	;
						10'd104	:	dt	<=	136	;
						10'd105	:	dt	<=	136	;
						10'd106	:	dt	<=	134	;
						10'd107	:	dt	<=	132	;
						10'd108	:	dt	<=	130	;
						10'd109	:	dt	<=	128	;
						10'd110	:	dt	<=	125	;
						10'd111	:	dt	<=	123	;
						10'd112	:	dt	<=	149	;
						10'd113	:	dt	<=	149	;
						10'd114	:	dt	<=	149	;
						10'd115	:	dt	<=	151	;
						10'd116	:	dt	<=	152	;
						10'd117	:	dt	<=	152	;
						10'd118	:	dt	<=	152	;
						10'd119	:	dt	<=	153	;
						10'd120	:	dt	<=	152	;
						10'd121	:	dt	<=	151	;
						10'd122	:	dt	<=	151	;
						10'd123	:	dt	<=	150	;
						10'd124	:	dt	<=	149	;
						10'd125	:	dt	<=	149	;
						10'd126	:	dt	<=	148	;
						10'd127	:	dt	<=	148	;
						10'd128	:	dt	<=	130	;
						10'd129	:	dt	<=	51	;
						10'd130	:	dt	<=	50	;
						10'd131	:	dt	<=	149	;
						10'd132	:	dt	<=	139	;
						10'd133	:	dt	<=	139	;
						10'd134	:	dt	<=	138	;
						10'd135	:	dt	<=	136	;
						10'd136	:	dt	<=	134	;
						10'd137	:	dt	<=	131	;
						10'd138	:	dt	<=	129	;
						10'd139	:	dt	<=	126	;
						10'd140	:	dt	<=	152	;
						10'd141	:	dt	<=	153	;
						10'd142	:	dt	<=	153	;
						10'd143	:	dt	<=	153	;
						10'd144	:	dt	<=	154	;
						10'd145	:	dt	<=	156	;
						10'd146	:	dt	<=	155	;
						10'd147	:	dt	<=	155	;
						10'd148	:	dt	<=	155	;
						10'd149	:	dt	<=	154	;
						10'd150	:	dt	<=	154	;
						10'd151	:	dt	<=	154	;
						10'd152	:	dt	<=	154	;
						10'd153	:	dt	<=	153	;
						10'd154	:	dt	<=	151	;
						10'd155	:	dt	<=	150	;
						10'd156	:	dt	<=	130	;
						10'd157	:	dt	<=	58	;
						10'd158	:	dt	<=	46	;
						10'd159	:	dt	<=	148	;
						10'd160	:	dt	<=	142	;
						10'd161	:	dt	<=	141	;
						10'd162	:	dt	<=	140	;
						10'd163	:	dt	<=	139	;
						10'd164	:	dt	<=	137	;
						10'd165	:	dt	<=	135	;
						10'd166	:	dt	<=	131	;
						10'd167	:	dt	<=	129	;
						10'd168	:	dt	<=	155	;
						10'd169	:	dt	<=	156	;
						10'd170	:	dt	<=	157	;
						10'd171	:	dt	<=	157	;
						10'd172	:	dt	<=	157	;
						10'd173	:	dt	<=	158	;
						10'd174	:	dt	<=	158	;
						10'd175	:	dt	<=	159	;
						10'd176	:	dt	<=	158	;
						10'd177	:	dt	<=	158	;
						10'd178	:	dt	<=	158	;
						10'd179	:	dt	<=	157	;
						10'd180	:	dt	<=	157	;
						10'd181	:	dt	<=	156	;
						10'd182	:	dt	<=	153	;
						10'd183	:	dt	<=	155	;
						10'd184	:	dt	<=	140	;
						10'd185	:	dt	<=	67	;
						10'd186	:	dt	<=	40	;
						10'd187	:	dt	<=	147	;
						10'd188	:	dt	<=	147	;
						10'd189	:	dt	<=	144	;
						10'd190	:	dt	<=	142	;
						10'd191	:	dt	<=	140	;
						10'd192	:	dt	<=	140	;
						10'd193	:	dt	<=	138	;
						10'd194	:	dt	<=	135	;
						10'd195	:	dt	<=	133	;
						10'd196	:	dt	<=	158	;
						10'd197	:	dt	<=	159	;
						10'd198	:	dt	<=	160	;
						10'd199	:	dt	<=	160	;
						10'd200	:	dt	<=	160	;
						10'd201	:	dt	<=	161	;
						10'd202	:	dt	<=	161	;
						10'd203	:	dt	<=	161	;
						10'd204	:	dt	<=	161	;
						10'd205	:	dt	<=	161	;
						10'd206	:	dt	<=	160	;
						10'd207	:	dt	<=	161	;
						10'd208	:	dt	<=	160	;
						10'd209	:	dt	<=	159	;
						10'd210	:	dt	<=	157	;
						10'd211	:	dt	<=	156	;
						10'd212	:	dt	<=	136	;
						10'd213	:	dt	<=	52	;
						10'd214	:	dt	<=	40	;
						10'd215	:	dt	<=	153	;
						10'd216	:	dt	<=	149	;
						10'd217	:	dt	<=	147	;
						10'd218	:	dt	<=	145	;
						10'd219	:	dt	<=	144	;
						10'd220	:	dt	<=	143	;
						10'd221	:	dt	<=	141	;
						10'd222	:	dt	<=	139	;
						10'd223	:	dt	<=	136	;
						10'd224	:	dt	<=	160	;
						10'd225	:	dt	<=	162	;
						10'd226	:	dt	<=	163	;
						10'd227	:	dt	<=	163	;
						10'd228	:	dt	<=	163	;
						10'd229	:	dt	<=	163	;
						10'd230	:	dt	<=	163	;
						10'd231	:	dt	<=	162	;
						10'd232	:	dt	<=	162	;
						10'd233	:	dt	<=	161	;
						10'd234	:	dt	<=	163	;
						10'd235	:	dt	<=	163	;
						10'd236	:	dt	<=	163	;
						10'd237	:	dt	<=	162	;
						10'd238	:	dt	<=	161	;
						10'd239	:	dt	<=	155	;
						10'd240	:	dt	<=	124	;
						10'd241	:	dt	<=	68	;
						10'd242	:	dt	<=	48	;
						10'd243	:	dt	<=	142	;
						10'd244	:	dt	<=	154	;
						10'd245	:	dt	<=	149	;
						10'd246	:	dt	<=	148	;
						10'd247	:	dt	<=	147	;
						10'd248	:	dt	<=	146	;
						10'd249	:	dt	<=	144	;
						10'd250	:	dt	<=	142	;
						10'd251	:	dt	<=	138	;
						10'd252	:	dt	<=	162	;
						10'd253	:	dt	<=	162	;
						10'd254	:	dt	<=	163	;
						10'd255	:	dt	<=	165	;
						10'd256	:	dt	<=	165	;
						10'd257	:	dt	<=	166	;
						10'd258	:	dt	<=	166	;
						10'd259	:	dt	<=	165	;
						10'd260	:	dt	<=	165	;
						10'd261	:	dt	<=	165	;
						10'd262	:	dt	<=	166	;
						10'd263	:	dt	<=	166	;
						10'd264	:	dt	<=	165	;
						10'd265	:	dt	<=	165	;
						10'd266	:	dt	<=	163	;
						10'd267	:	dt	<=	158	;
						10'd268	:	dt	<=	138	;
						10'd269	:	dt	<=	98	;
						10'd270	:	dt	<=	43	;
						10'd271	:	dt	<=	125	;
						10'd272	:	dt	<=	161	;
						10'd273	:	dt	<=	152	;
						10'd274	:	dt	<=	152	;
						10'd275	:	dt	<=	150	;
						10'd276	:	dt	<=	148	;
						10'd277	:	dt	<=	147	;
						10'd278	:	dt	<=	143	;
						10'd279	:	dt	<=	140	;
						10'd280	:	dt	<=	163	;
						10'd281	:	dt	<=	165	;
						10'd282	:	dt	<=	165	;
						10'd283	:	dt	<=	166	;
						10'd284	:	dt	<=	166	;
						10'd285	:	dt	<=	168	;
						10'd286	:	dt	<=	168	;
						10'd287	:	dt	<=	168	;
						10'd288	:	dt	<=	168	;
						10'd289	:	dt	<=	168	;
						10'd290	:	dt	<=	169	;
						10'd291	:	dt	<=	168	;
						10'd292	:	dt	<=	167	;
						10'd293	:	dt	<=	166	;
						10'd294	:	dt	<=	166	;
						10'd295	:	dt	<=	159	;
						10'd296	:	dt	<=	142	;
						10'd297	:	dt	<=	96	;
						10'd298	:	dt	<=	30	;
						10'd299	:	dt	<=	112	;
						10'd300	:	dt	<=	166	;
						10'd301	:	dt	<=	152	;
						10'd302	:	dt	<=	153	;
						10'd303	:	dt	<=	153	;
						10'd304	:	dt	<=	150	;
						10'd305	:	dt	<=	148	;
						10'd306	:	dt	<=	146	;
						10'd307	:	dt	<=	142	;
						10'd308	:	dt	<=	166	;
						10'd309	:	dt	<=	166	;
						10'd310	:	dt	<=	167	;
						10'd311	:	dt	<=	167	;
						10'd312	:	dt	<=	167	;
						10'd313	:	dt	<=	168	;
						10'd314	:	dt	<=	170	;
						10'd315	:	dt	<=	169	;
						10'd316	:	dt	<=	169	;
						10'd317	:	dt	<=	169	;
						10'd318	:	dt	<=	169	;
						10'd319	:	dt	<=	170	;
						10'd320	:	dt	<=	168	;
						10'd321	:	dt	<=	169	;
						10'd322	:	dt	<=	167	;
						10'd323	:	dt	<=	163	;
						10'd324	:	dt	<=	153	;
						10'd325	:	dt	<=	97	;
						10'd326	:	dt	<=	34	;
						10'd327	:	dt	<=	83	;
						10'd328	:	dt	<=	173	;
						10'd329	:	dt	<=	152	;
						10'd330	:	dt	<=	155	;
						10'd331	:	dt	<=	154	;
						10'd332	:	dt	<=	152	;
						10'd333	:	dt	<=	150	;
						10'd334	:	dt	<=	148	;
						10'd335	:	dt	<=	145	;
						10'd336	:	dt	<=	168	;
						10'd337	:	dt	<=	168	;
						10'd338	:	dt	<=	169	;
						10'd339	:	dt	<=	169	;
						10'd340	:	dt	<=	168	;
						10'd341	:	dt	<=	169	;
						10'd342	:	dt	<=	170	;
						10'd343	:	dt	<=	171	;
						10'd344	:	dt	<=	171	;
						10'd345	:	dt	<=	170	;
						10'd346	:	dt	<=	171	;
						10'd347	:	dt	<=	172	;
						10'd348	:	dt	<=	173	;
						10'd349	:	dt	<=	165	;
						10'd350	:	dt	<=	147	;
						10'd351	:	dt	<=	134	;
						10'd352	:	dt	<=	127	;
						10'd353	:	dt	<=	124	;
						10'd354	:	dt	<=	73	;
						10'd355	:	dt	<=	103	;
						10'd356	:	dt	<=	147	;
						10'd357	:	dt	<=	167	;
						10'd358	:	dt	<=	156	;
						10'd359	:	dt	<=	155	;
						10'd360	:	dt	<=	153	;
						10'd361	:	dt	<=	151	;
						10'd362	:	dt	<=	149	;
						10'd363	:	dt	<=	146	;
						10'd364	:	dt	<=	169	;
						10'd365	:	dt	<=	169	;
						10'd366	:	dt	<=	169	;
						10'd367	:	dt	<=	170	;
						10'd368	:	dt	<=	171	;
						10'd369	:	dt	<=	171	;
						10'd370	:	dt	<=	172	;
						10'd371	:	dt	<=	173	;
						10'd372	:	dt	<=	173	;
						10'd373	:	dt	<=	172	;
						10'd374	:	dt	<=	175	;
						10'd375	:	dt	<=	174	;
						10'd376	:	dt	<=	165	;
						10'd377	:	dt	<=	156	;
						10'd378	:	dt	<=	147	;
						10'd379	:	dt	<=	94	;
						10'd380	:	dt	<=	48	;
						10'd381	:	dt	<=	106	;
						10'd382	:	dt	<=	118	;
						10'd383	:	dt	<=	149	;
						10'd384	:	dt	<=	72	;
						10'd385	:	dt	<=	132	;
						10'd386	:	dt	<=	167	;
						10'd387	:	dt	<=	157	;
						10'd388	:	dt	<=	156	;
						10'd389	:	dt	<=	154	;
						10'd390	:	dt	<=	151	;
						10'd391	:	dt	<=	148	;
						10'd392	:	dt	<=	170	;
						10'd393	:	dt	<=	170	;
						10'd394	:	dt	<=	171	;
						10'd395	:	dt	<=	172	;
						10'd396	:	dt	<=	173	;
						10'd397	:	dt	<=	173	;
						10'd398	:	dt	<=	174	;
						10'd399	:	dt	<=	173	;
						10'd400	:	dt	<=	174	;
						10'd401	:	dt	<=	176	;
						10'd402	:	dt	<=	168	;
						10'd403	:	dt	<=	149	;
						10'd404	:	dt	<=	97	;
						10'd405	:	dt	<=	111	;
						10'd406	:	dt	<=	149	;
						10'd407	:	dt	<=	93	;
						10'd408	:	dt	<=	44	;
						10'd409	:	dt	<=	59	;
						10'd410	:	dt	<=	121	;
						10'd411	:	dt	<=	120	;
						10'd412	:	dt	<=	44	;
						10'd413	:	dt	<=	16	;
						10'd414	:	dt	<=	102	;
						10'd415	:	dt	<=	167	;
						10'd416	:	dt	<=	156	;
						10'd417	:	dt	<=	155	;
						10'd418	:	dt	<=	153	;
						10'd419	:	dt	<=	150	;
						10'd420	:	dt	<=	172	;
						10'd421	:	dt	<=	172	;
						10'd422	:	dt	<=	173	;
						10'd423	:	dt	<=	174	;
						10'd424	:	dt	<=	175	;
						10'd425	:	dt	<=	176	;
						10'd426	:	dt	<=	175	;
						10'd427	:	dt	<=	175	;
						10'd428	:	dt	<=	177	;
						10'd429	:	dt	<=	168	;
						10'd430	:	dt	<=	157	;
						10'd431	:	dt	<=	140	;
						10'd432	:	dt	<=	87	;
						10'd433	:	dt	<=	56	;
						10'd434	:	dt	<=	109	;
						10'd435	:	dt	<=	122	;
						10'd436	:	dt	<=	70	;
						10'd437	:	dt	<=	39	;
						10'd438	:	dt	<=	93	;
						10'd439	:	dt	<=	102	;
						10'd440	:	dt	<=	52	;
						10'd441	:	dt	<=	21	;
						10'd442	:	dt	<=	25	;
						10'd443	:	dt	<=	153	;
						10'd444	:	dt	<=	162	;
						10'd445	:	dt	<=	156	;
						10'd446	:	dt	<=	154	;
						10'd447	:	dt	<=	153	;
						10'd448	:	dt	<=	173	;
						10'd449	:	dt	<=	173	;
						10'd450	:	dt	<=	174	;
						10'd451	:	dt	<=	175	;
						10'd452	:	dt	<=	176	;
						10'd453	:	dt	<=	176	;
						10'd454	:	dt	<=	175	;
						10'd455	:	dt	<=	177	;
						10'd456	:	dt	<=	175	;
						10'd457	:	dt	<=	159	;
						10'd458	:	dt	<=	143	;
						10'd459	:	dt	<=	117	;
						10'd460	:	dt	<=	112	;
						10'd461	:	dt	<=	90	;
						10'd462	:	dt	<=	70	;
						10'd463	:	dt	<=	130	;
						10'd464	:	dt	<=	83	;
						10'd465	:	dt	<=	31	;
						10'd466	:	dt	<=	36	;
						10'd467	:	dt	<=	65	;
						10'd468	:	dt	<=	68	;
						10'd469	:	dt	<=	30	;
						10'd470	:	dt	<=	19	;
						10'd471	:	dt	<=	140	;
						10'd472	:	dt	<=	167	;
						10'd473	:	dt	<=	157	;
						10'd474	:	dt	<=	157	;
						10'd475	:	dt	<=	154	;
						10'd476	:	dt	<=	174	;
						10'd477	:	dt	<=	174	;
						10'd478	:	dt	<=	174	;
						10'd479	:	dt	<=	175	;
						10'd480	:	dt	<=	176	;
						10'd481	:	dt	<=	176	;
						10'd482	:	dt	<=	176	;
						10'd483	:	dt	<=	178	;
						10'd484	:	dt	<=	171	;
						10'd485	:	dt	<=	150	;
						10'd486	:	dt	<=	114	;
						10'd487	:	dt	<=	71	;
						10'd488	:	dt	<=	95	;
						10'd489	:	dt	<=	97	;
						10'd490	:	dt	<=	52	;
						10'd491	:	dt	<=	92	;
						10'd492	:	dt	<=	97	;
						10'd493	:	dt	<=	36	;
						10'd494	:	dt	<=	24	;
						10'd495	:	dt	<=	46	;
						10'd496	:	dt	<=	86	;
						10'd497	:	dt	<=	44	;
						10'd498	:	dt	<=	11	;
						10'd499	:	dt	<=	129	;
						10'd500	:	dt	<=	170	;
						10'd501	:	dt	<=	158	;
						10'd502	:	dt	<=	157	;
						10'd503	:	dt	<=	155	;
						10'd504	:	dt	<=	173	;
						10'd505	:	dt	<=	174	;
						10'd506	:	dt	<=	174	;
						10'd507	:	dt	<=	175	;
						10'd508	:	dt	<=	177	;
						10'd509	:	dt	<=	178	;
						10'd510	:	dt	<=	179	;
						10'd511	:	dt	<=	180	;
						10'd512	:	dt	<=	175	;
						10'd513	:	dt	<=	149	;
						10'd514	:	dt	<=	131	;
						10'd515	:	dt	<=	69	;
						10'd516	:	dt	<=	34	;
						10'd517	:	dt	<=	74	;
						10'd518	:	dt	<=	14	;
						10'd519	:	dt	<=	48	;
						10'd520	:	dt	<=	91	;
						10'd521	:	dt	<=	23	;
						10'd522	:	dt	<=	28	;
						10'd523	:	dt	<=	43	;
						10'd524	:	dt	<=	93	;
						10'd525	:	dt	<=	80	;
						10'd526	:	dt	<=	13	;
						10'd527	:	dt	<=	104	;
						10'd528	:	dt	<=	174	;
						10'd529	:	dt	<=	159	;
						10'd530	:	dt	<=	159	;
						10'd531	:	dt	<=	157	;
						10'd532	:	dt	<=	173	;
						10'd533	:	dt	<=	174	;
						10'd534	:	dt	<=	174	;
						10'd535	:	dt	<=	176	;
						10'd536	:	dt	<=	177	;
						10'd537	:	dt	<=	178	;
						10'd538	:	dt	<=	180	;
						10'd539	:	dt	<=	179	;
						10'd540	:	dt	<=	182	;
						10'd541	:	dt	<=	153	;
						10'd542	:	dt	<=	121	;
						10'd543	:	dt	<=	92	;
						10'd544	:	dt	<=	59	;
						10'd545	:	dt	<=	38	;
						10'd546	:	dt	<=	15	;
						10'd547	:	dt	<=	43	;
						10'd548	:	dt	<=	51	;
						10'd549	:	dt	<=	6	;
						10'd550	:	dt	<=	37	;
						10'd551	:	dt	<=	87	;
						10'd552	:	dt	<=	109	;
						10'd553	:	dt	<=	96	;
						10'd554	:	dt	<=	19	;
						10'd555	:	dt	<=	107	;
						10'd556	:	dt	<=	175	;
						10'd557	:	dt	<=	160	;
						10'd558	:	dt	<=	161	;
						10'd559	:	dt	<=	158	;
						10'd560	:	dt	<=	173	;
						10'd561	:	dt	<=	174	;
						10'd562	:	dt	<=	175	;
						10'd563	:	dt	<=	175	;
						10'd564	:	dt	<=	176	;
						10'd565	:	dt	<=	177	;
						10'd566	:	dt	<=	178	;
						10'd567	:	dt	<=	179	;
						10'd568	:	dt	<=	184	;
						10'd569	:	dt	<=	153	;
						10'd570	:	dt	<=	132	;
						10'd571	:	dt	<=	126	;
						10'd572	:	dt	<=	88	;
						10'd573	:	dt	<=	46	;
						10'd574	:	dt	<=	46	;
						10'd575	:	dt	<=	68	;
						10'd576	:	dt	<=	57	;
						10'd577	:	dt	<=	45	;
						10'd578	:	dt	<=	117	;
						10'd579	:	dt	<=	126	;
						10'd580	:	dt	<=	109	;
						10'd581	:	dt	<=	60	;
						10'd582	:	dt	<=	39	;
						10'd583	:	dt	<=	161	;
						10'd584	:	dt	<=	165	;
						10'd585	:	dt	<=	161	;
						10'd586	:	dt	<=	159	;
						10'd587	:	dt	<=	155	;
						10'd588	:	dt	<=	174	;
						10'd589	:	dt	<=	175	;
						10'd590	:	dt	<=	176	;
						10'd591	:	dt	<=	176	;
						10'd592	:	dt	<=	178	;
						10'd593	:	dt	<=	179	;
						10'd594	:	dt	<=	179	;
						10'd595	:	dt	<=	179	;
						10'd596	:	dt	<=	183	;
						10'd597	:	dt	<=	161	;
						10'd598	:	dt	<=	125	;
						10'd599	:	dt	<=	126	;
						10'd600	:	dt	<=	100	;
						10'd601	:	dt	<=	68	;
						10'd602	:	dt	<=	58	;
						10'd603	:	dt	<=	83	;
						10'd604	:	dt	<=	132	;
						10'd605	:	dt	<=	139	;
						10'd606	:	dt	<=	148	;
						10'd607	:	dt	<=	111	;
						10'd608	:	dt	<=	79	;
						10'd609	:	dt	<=	23	;
						10'd610	:	dt	<=	101	;
						10'd611	:	dt	<=	177	;
						10'd612	:	dt	<=	157	;
						10'd613	:	dt	<=	159	;
						10'd614	:	dt	<=	162	;
						10'd615	:	dt	<=	164	;
						10'd616	:	dt	<=	173	;
						10'd617	:	dt	<=	173	;
						10'd618	:	dt	<=	174	;
						10'd619	:	dt	<=	176	;
						10'd620	:	dt	<=	177	;
						10'd621	:	dt	<=	178	;
						10'd622	:	dt	<=	179	;
						10'd623	:	dt	<=	178	;
						10'd624	:	dt	<=	183	;
						10'd625	:	dt	<=	171	;
						10'd626	:	dt	<=	122	;
						10'd627	:	dt	<=	123	;
						10'd628	:	dt	<=	104	;
						10'd629	:	dt	<=	75	;
						10'd630	:	dt	<=	61	;
						10'd631	:	dt	<=	69	;
						10'd632	:	dt	<=	139	;
						10'd633	:	dt	<=	137	;
						10'd634	:	dt	<=	120	;
						10'd635	:	dt	<=	87	;
						10'd636	:	dt	<=	46	;
						10'd637	:	dt	<=	22	;
						10'd638	:	dt	<=	149	;
						10'd639	:	dt	<=	173	;
						10'd640	:	dt	<=	171	;
						10'd641	:	dt	<=	171	;
						10'd642	:	dt	<=	149	;
						10'd643	:	dt	<=	110	;
						10'd644	:	dt	<=	180	;
						10'd645	:	dt	<=	180	;
						10'd646	:	dt	<=	181	;
						10'd647	:	dt	<=	181	;
						10'd648	:	dt	<=	182	;
						10'd649	:	dt	<=	183	;
						10'd650	:	dt	<=	184	;
						10'd651	:	dt	<=	184	;
						10'd652	:	dt	<=	184	;
						10'd653	:	dt	<=	187	;
						10'd654	:	dt	<=	131	;
						10'd655	:	dt	<=	101	;
						10'd656	:	dt	<=	96	;
						10'd657	:	dt	<=	75	;
						10'd658	:	dt	<=	67	;
						10'd659	:	dt	<=	64	;
						10'd660	:	dt	<=	118	;
						10'd661	:	dt	<=	120	;
						10'd662	:	dt	<=	98	;
						10'd663	:	dt	<=	63	;
						10'd664	:	dt	<=	15	;
						10'd665	:	dt	<=	82	;
						10'd666	:	dt	<=	182	;
						10'd667	:	dt	<=	150	;
						10'd668	:	dt	<=	125	;
						10'd669	:	dt	<=	87	;
						10'd670	:	dt	<=	36	;
						10'd671	:	dt	<=	13	;
						10'd672	:	dt	<=	134	;
						10'd673	:	dt	<=	139	;
						10'd674	:	dt	<=	144	;
						10'd675	:	dt	<=	147	;
						10'd676	:	dt	<=	153	;
						10'd677	:	dt	<=	158	;
						10'd678	:	dt	<=	162	;
						10'd679	:	dt	<=	165	;
						10'd680	:	dt	<=	167	;
						10'd681	:	dt	<=	174	;
						10'd682	:	dt	<=	157	;
						10'd683	:	dt	<=	96	;
						10'd684	:	dt	<=	94	;
						10'd685	:	dt	<=	86	;
						10'd686	:	dt	<=	82	;
						10'd687	:	dt	<=	60	;
						10'd688	:	dt	<=	87	;
						10'd689	:	dt	<=	100	;
						10'd690	:	dt	<=	75	;
						10'd691	:	dt	<=	29	;
						10'd692	:	dt	<=	37	;
						10'd693	:	dt	<=	115	;
						10'd694	:	dt	<=	68	;
						10'd695	:	dt	<=	32	;
						10'd696	:	dt	<=	10	;
						10'd697	:	dt	<=	2	;
						10'd698	:	dt	<=	2	;
						10'd699	:	dt	<=	8	;
						10'd700	:	dt	<=	61	;
						10'd701	:	dt	<=	62	;
						10'd702	:	dt	<=	64	;
						10'd703	:	dt	<=	64	;
						10'd704	:	dt	<=	65	;
						10'd705	:	dt	<=	69	;
						10'd706	:	dt	<=	69	;
						10'd707	:	dt	<=	70	;
						10'd708	:	dt	<=	70	;
						10'd709	:	dt	<=	69	;
						10'd710	:	dt	<=	83	;
						10'd711	:	dt	<=	119	;
						10'd712	:	dt	<=	94	;
						10'd713	:	dt	<=	91	;
						10'd714	:	dt	<=	75	;
						10'd715	:	dt	<=	50	;
						10'd716	:	dt	<=	50	;
						10'd717	:	dt	<=	50	;
						10'd718	:	dt	<=	25	;
						10'd719	:	dt	<=	11	;
						10'd720	:	dt	<=	37	;
						10'd721	:	dt	<=	24	;
						10'd722	:	dt	<=	3	;
						10'd723	:	dt	<=	0	;
						10'd724	:	dt	<=	6	;
						10'd725	:	dt	<=	0	;
						10'd726	:	dt	<=	0	;
						10'd727	:	dt	<=	0	;
						10'd728	:	dt	<=	71	;
						10'd729	:	dt	<=	70	;
						10'd730	:	dt	<=	71	;
						10'd731	:	dt	<=	72	;
						10'd732	:	dt	<=	70	;
						10'd733	:	dt	<=	70	;
						10'd734	:	dt	<=	77	;
						10'd735	:	dt	<=	74	;
						10'd736	:	dt	<=	75	;
						10'd737	:	dt	<=	70	;
						10'd738	:	dt	<=	92	;
						10'd739	:	dt	<=	144	;
						10'd740	:	dt	<=	123	;
						10'd741	:	dt	<=	94	;
						10'd742	:	dt	<=	61	;
						10'd743	:	dt	<=	45	;
						10'd744	:	dt	<=	44	;
						10'd745	:	dt	<=	42	;
						10'd746	:	dt	<=	18	;
						10'd747	:	dt	<=	18	;
						10'd748	:	dt	<=	20	;
						10'd749	:	dt	<=	11	;
						10'd750	:	dt	<=	14	;
						10'd751	:	dt	<=	0	;
						10'd752	:	dt	<=	0	;
						10'd753	:	dt	<=	0	;
						10'd754	:	dt	<=	0	;
						10'd755	:	dt	<=	0	;
						10'd756	:	dt	<=	70	;
						10'd757	:	dt	<=	71	;
						10'd758	:	dt	<=	71	;
						10'd759	:	dt	<=	72	;
						10'd760	:	dt	<=	72	;
						10'd761	:	dt	<=	72	;
						10'd762	:	dt	<=	80	;
						10'd763	:	dt	<=	77	;
						10'd764	:	dt	<=	80	;
						10'd765	:	dt	<=	75	;
						10'd766	:	dt	<=	110	;
						10'd767	:	dt	<=	130	;
						10'd768	:	dt	<=	128	;
						10'd769	:	dt	<=	102	;
						10'd770	:	dt	<=	78	;
						10'd771	:	dt	<=	66	;
						10'd772	:	dt	<=	53	;
						10'd773	:	dt	<=	40	;
						10'd774	:	dt	<=	14	;
						10'd775	:	dt	<=	16	;
						10'd776	:	dt	<=	12	;
						10'd777	:	dt	<=	8	;
						10'd778	:	dt	<=	2	;
						10'd779	:	dt	<=	2	;
						10'd780	:	dt	<=	0	;
						10'd781	:	dt	<=	0	;
						10'd782	:	dt	<=	0	;
						10'd783	:	dt	<=	0	;
					endcase
				end
				2'd2	:	begin
					case (cnt)
						10'd0	:	dt	<=	125	;
						10'd1	:	dt	<=	126	;
						10'd2	:	dt	<=	132	;
						10'd3	:	dt	<=	138	;
						10'd4	:	dt	<=	142	;
						10'd5	:	dt	<=	144	;
						10'd6	:	dt	<=	148	;
						10'd7	:	dt	<=	151	;
						10'd8	:	dt	<=	153	;
						10'd9	:	dt	<=	154	;
						10'd10	:	dt	<=	156	;
						10'd11	:	dt	<=	157	;
						10'd12	:	dt	<=	159	;
						10'd13	:	dt	<=	160	;
						10'd14	:	dt	<=	161	;
						10'd15	:	dt	<=	161	;
						10'd16	:	dt	<=	162	;
						10'd17	:	dt	<=	162	;
						10'd18	:	dt	<=	161	;
						10'd19	:	dt	<=	162	;
						10'd20	:	dt	<=	162	;
						10'd21	:	dt	<=	161	;
						10'd22	:	dt	<=	162	;
						10'd23	:	dt	<=	161	;
						10'd24	:	dt	<=	160	;
						10'd25	:	dt	<=	159	;
						10'd26	:	dt	<=	157	;
						10'd27	:	dt	<=	158	;
						10'd28	:	dt	<=	126	;
						10'd29	:	dt	<=	127	;
						10'd30	:	dt	<=	133	;
						10'd31	:	dt	<=	138	;
						10'd32	:	dt	<=	143	;
						10'd33	:	dt	<=	145	;
						10'd34	:	dt	<=	148	;
						10'd35	:	dt	<=	151	;
						10'd36	:	dt	<=	153	;
						10'd37	:	dt	<=	155	;
						10'd38	:	dt	<=	157	;
						10'd39	:	dt	<=	158	;
						10'd40	:	dt	<=	160	;
						10'd41	:	dt	<=	161	;
						10'd42	:	dt	<=	161	;
						10'd43	:	dt	<=	162	;
						10'd44	:	dt	<=	162	;
						10'd45	:	dt	<=	162	;
						10'd46	:	dt	<=	162	;
						10'd47	:	dt	<=	163	;
						10'd48	:	dt	<=	164	;
						10'd49	:	dt	<=	163	;
						10'd50	:	dt	<=	162	;
						10'd51	:	dt	<=	162	;
						10'd52	:	dt	<=	161	;
						10'd53	:	dt	<=	161	;
						10'd54	:	dt	<=	158	;
						10'd55	:	dt	<=	158	;
						10'd56	:	dt	<=	127	;
						10'd57	:	dt	<=	128	;
						10'd58	:	dt	<=	134	;
						10'd59	:	dt	<=	139	;
						10'd60	:	dt	<=	144	;
						10'd61	:	dt	<=	147	;
						10'd62	:	dt	<=	149	;
						10'd63	:	dt	<=	152	;
						10'd64	:	dt	<=	155	;
						10'd65	:	dt	<=	156	;
						10'd66	:	dt	<=	159	;
						10'd67	:	dt	<=	159	;
						10'd68	:	dt	<=	161	;
						10'd69	:	dt	<=	162	;
						10'd70	:	dt	<=	163	;
						10'd71	:	dt	<=	162	;
						10'd72	:	dt	<=	164	;
						10'd73	:	dt	<=	163	;
						10'd74	:	dt	<=	164	;
						10'd75	:	dt	<=	165	;
						10'd76	:	dt	<=	166	;
						10'd77	:	dt	<=	165	;
						10'd78	:	dt	<=	164	;
						10'd79	:	dt	<=	163	;
						10'd80	:	dt	<=	163	;
						10'd81	:	dt	<=	161	;
						10'd82	:	dt	<=	160	;
						10'd83	:	dt	<=	160	;
						10'd84	:	dt	<=	127	;
						10'd85	:	dt	<=	129	;
						10'd86	:	dt	<=	136	;
						10'd87	:	dt	<=	140	;
						10'd88	:	dt	<=	144	;
						10'd89	:	dt	<=	147	;
						10'd90	:	dt	<=	150	;
						10'd91	:	dt	<=	154	;
						10'd92	:	dt	<=	155	;
						10'd93	:	dt	<=	158	;
						10'd94	:	dt	<=	161	;
						10'd95	:	dt	<=	159	;
						10'd96	:	dt	<=	161	;
						10'd97	:	dt	<=	160	;
						10'd98	:	dt	<=	162	;
						10'd99	:	dt	<=	166	;
						10'd100	:	dt	<=	164	;
						10'd101	:	dt	<=	165	;
						10'd102	:	dt	<=	165	;
						10'd103	:	dt	<=	166	;
						10'd104	:	dt	<=	166	;
						10'd105	:	dt	<=	165	;
						10'd106	:	dt	<=	164	;
						10'd107	:	dt	<=	164	;
						10'd108	:	dt	<=	163	;
						10'd109	:	dt	<=	162	;
						10'd110	:	dt	<=	162	;
						10'd111	:	dt	<=	162	;
						10'd112	:	dt	<=	127	;
						10'd113	:	dt	<=	130	;
						10'd114	:	dt	<=	136	;
						10'd115	:	dt	<=	142	;
						10'd116	:	dt	<=	146	;
						10'd117	:	dt	<=	149	;
						10'd118	:	dt	<=	152	;
						10'd119	:	dt	<=	155	;
						10'd120	:	dt	<=	157	;
						10'd121	:	dt	<=	158	;
						10'd122	:	dt	<=	160	;
						10'd123	:	dt	<=	161	;
						10'd124	:	dt	<=	193	;
						10'd125	:	dt	<=	175	;
						10'd126	:	dt	<=	128	;
						10'd127	:	dt	<=	152	;
						10'd128	:	dt	<=	169	;
						10'd129	:	dt	<=	164	;
						10'd130	:	dt	<=	167	;
						10'd131	:	dt	<=	169	;
						10'd132	:	dt	<=	166	;
						10'd133	:	dt	<=	166	;
						10'd134	:	dt	<=	166	;
						10'd135	:	dt	<=	165	;
						10'd136	:	dt	<=	165	;
						10'd137	:	dt	<=	164	;
						10'd138	:	dt	<=	163	;
						10'd139	:	dt	<=	162	;
						10'd140	:	dt	<=	128	;
						10'd141	:	dt	<=	130	;
						10'd142	:	dt	<=	136	;
						10'd143	:	dt	<=	142	;
						10'd144	:	dt	<=	147	;
						10'd145	:	dt	<=	150	;
						10'd146	:	dt	<=	152	;
						10'd147	:	dt	<=	155	;
						10'd148	:	dt	<=	157	;
						10'd149	:	dt	<=	157	;
						10'd150	:	dt	<=	158	;
						10'd151	:	dt	<=	171	;
						10'd152	:	dt	<=	223	;
						10'd153	:	dt	<=	202	;
						10'd154	:	dt	<=	145	;
						10'd155	:	dt	<=	123	;
						10'd156	:	dt	<=	174	;
						10'd157	:	dt	<=	170	;
						10'd158	:	dt	<=	147	;
						10'd159	:	dt	<=	148	;
						10'd160	:	dt	<=	170	;
						10'd161	:	dt	<=	166	;
						10'd162	:	dt	<=	167	;
						10'd163	:	dt	<=	167	;
						10'd164	:	dt	<=	167	;
						10'd165	:	dt	<=	165	;
						10'd166	:	dt	<=	163	;
						10'd167	:	dt	<=	163	;
						10'd168	:	dt	<=	128	;
						10'd169	:	dt	<=	132	;
						10'd170	:	dt	<=	136	;
						10'd171	:	dt	<=	142	;
						10'd172	:	dt	<=	147	;
						10'd173	:	dt	<=	151	;
						10'd174	:	dt	<=	154	;
						10'd175	:	dt	<=	156	;
						10'd176	:	dt	<=	154	;
						10'd177	:	dt	<=	167	;
						10'd178	:	dt	<=	163	;
						10'd179	:	dt	<=	158	;
						10'd180	:	dt	<=	217	;
						10'd181	:	dt	<=	206	;
						10'd182	:	dt	<=	168	;
						10'd183	:	dt	<=	121	;
						10'd184	:	dt	<=	138	;
						10'd185	:	dt	<=	155	;
						10'd186	:	dt	<=	127	;
						10'd187	:	dt	<=	87	;
						10'd188	:	dt	<=	153	;
						10'd189	:	dt	<=	172	;
						10'd190	:	dt	<=	167	;
						10'd191	:	dt	<=	168	;
						10'd192	:	dt	<=	167	;
						10'd193	:	dt	<=	166	;
						10'd194	:	dt	<=	165	;
						10'd195	:	dt	<=	164	;
						10'd196	:	dt	<=	128	;
						10'd197	:	dt	<=	132	;
						10'd198	:	dt	<=	137	;
						10'd199	:	dt	<=	141	;
						10'd200	:	dt	<=	147	;
						10'd201	:	dt	<=	152	;
						10'd202	:	dt	<=	154	;
						10'd203	:	dt	<=	151	;
						10'd204	:	dt	<=	172	;
						10'd205	:	dt	<=	206	;
						10'd206	:	dt	<=	164	;
						10'd207	:	dt	<=	134	;
						10'd208	:	dt	<=	172	;
						10'd209	:	dt	<=	179	;
						10'd210	:	dt	<=	153	;
						10'd211	:	dt	<=	92	;
						10'd212	:	dt	<=	121	;
						10'd213	:	dt	<=	118	;
						10'd214	:	dt	<=	96	;
						10'd215	:	dt	<=	74	;
						10'd216	:	dt	<=	120	;
						10'd217	:	dt	<=	177	;
						10'd218	:	dt	<=	166	;
						10'd219	:	dt	<=	168	;
						10'd220	:	dt	<=	167	;
						10'd221	:	dt	<=	167	;
						10'd222	:	dt	<=	167	;
						10'd223	:	dt	<=	166	;
						10'd224	:	dt	<=	129	;
						10'd225	:	dt	<=	132	;
						10'd226	:	dt	<=	138	;
						10'd227	:	dt	<=	143	;
						10'd228	:	dt	<=	148	;
						10'd229	:	dt	<=	149	;
						10'd230	:	dt	<=	167	;
						10'd231	:	dt	<=	153	;
						10'd232	:	dt	<=	178	;
						10'd233	:	dt	<=	213	;
						10'd234	:	dt	<=	176	;
						10'd235	:	dt	<=	130	;
						10'd236	:	dt	<=	149	;
						10'd237	:	dt	<=	168	;
						10'd238	:	dt	<=	137	;
						10'd239	:	dt	<=	90	;
						10'd240	:	dt	<=	131	;
						10'd241	:	dt	<=	103	;
						10'd242	:	dt	<=	77	;
						10'd243	:	dt	<=	71	;
						10'd244	:	dt	<=	115	;
						10'd245	:	dt	<=	178	;
						10'd246	:	dt	<=	167	;
						10'd247	:	dt	<=	169	;
						10'd248	:	dt	<=	169	;
						10'd249	:	dt	<=	168	;
						10'd250	:	dt	<=	168	;
						10'd251	:	dt	<=	167	;
						10'd252	:	dt	<=	130	;
						10'd253	:	dt	<=	134	;
						10'd254	:	dt	<=	140	;
						10'd255	:	dt	<=	145	;
						10'd256	:	dt	<=	146	;
						10'd257	:	dt	<=	159	;
						10'd258	:	dt	<=	210	;
						10'd259	:	dt	<=	159	;
						10'd260	:	dt	<=	126	;
						10'd261	:	dt	<=	195	;
						10'd262	:	dt	<=	194	;
						10'd263	:	dt	<=	145	;
						10'd264	:	dt	<=	116	;
						10'd265	:	dt	<=	174	;
						10'd266	:	dt	<=	173	;
						10'd267	:	dt	<=	159	;
						10'd268	:	dt	<=	148	;
						10'd269	:	dt	<=	121	;
						10'd270	:	dt	<=	74	;
						10'd271	:	dt	<=	57	;
						10'd272	:	dt	<=	120	;
						10'd273	:	dt	<=	179	;
						10'd274	:	dt	<=	170	;
						10'd275	:	dt	<=	169	;
						10'd276	:	dt	<=	169	;
						10'd277	:	dt	<=	168	;
						10'd278	:	dt	<=	168	;
						10'd279	:	dt	<=	167	;
						10'd280	:	dt	<=	131	;
						10'd281	:	dt	<=	135	;
						10'd282	:	dt	<=	141	;
						10'd283	:	dt	<=	147	;
						10'd284	:	dt	<=	141	;
						10'd285	:	dt	<=	186	;
						10'd286	:	dt	<=	213	;
						10'd287	:	dt	<=	174	;
						10'd288	:	dt	<=	128	;
						10'd289	:	dt	<=	152	;
						10'd290	:	dt	<=	200	;
						10'd291	:	dt	<=	156	;
						10'd292	:	dt	<=	92	;
						10'd293	:	dt	<=	101	;
						10'd294	:	dt	<=	168	;
						10'd295	:	dt	<=	173	;
						10'd296	:	dt	<=	158	;
						10'd297	:	dt	<=	159	;
						10'd298	:	dt	<=	128	;
						10'd299	:	dt	<=	61	;
						10'd300	:	dt	<=	134	;
						10'd301	:	dt	<=	179	;
						10'd302	:	dt	<=	171	;
						10'd303	:	dt	<=	170	;
						10'd304	:	dt	<=	170	;
						10'd305	:	dt	<=	169	;
						10'd306	:	dt	<=	168	;
						10'd307	:	dt	<=	168	;
						10'd308	:	dt	<=	132	;
						10'd309	:	dt	<=	134	;
						10'd310	:	dt	<=	140	;
						10'd311	:	dt	<=	146	;
						10'd312	:	dt	<=	147	;
						10'd313	:	dt	<=	190	;
						10'd314	:	dt	<=	196	;
						10'd315	:	dt	<=	187	;
						10'd316	:	dt	<=	143	;
						10'd317	:	dt	<=	113	;
						10'd318	:	dt	<=	188	;
						10'd319	:	dt	<=	160	;
						10'd320	:	dt	<=	114	;
						10'd321	:	dt	<=	41	;
						10'd322	:	dt	<=	90	;
						10'd323	:	dt	<=	127	;
						10'd324	:	dt	<=	154	;
						10'd325	:	dt	<=	172	;
						10'd326	:	dt	<=	174	;
						10'd327	:	dt	<=	114	;
						10'd328	:	dt	<=	141	;
						10'd329	:	dt	<=	180	;
						10'd330	:	dt	<=	171	;
						10'd331	:	dt	<=	172	;
						10'd332	:	dt	<=	172	;
						10'd333	:	dt	<=	171	;
						10'd334	:	dt	<=	170	;
						10'd335	:	dt	<=	168	;
						10'd336	:	dt	<=	130	;
						10'd337	:	dt	<=	133	;
						10'd338	:	dt	<=	138	;
						10'd339	:	dt	<=	142	;
						10'd340	:	dt	<=	150	;
						10'd341	:	dt	<=	194	;
						10'd342	:	dt	<=	180	;
						10'd343	:	dt	<=	184	;
						10'd344	:	dt	<=	152	;
						10'd345	:	dt	<=	100	;
						10'd346	:	dt	<=	154	;
						10'd347	:	dt	<=	178	;
						10'd348	:	dt	<=	124	;
						10'd349	:	dt	<=	54	;
						10'd350	:	dt	<=	50	;
						10'd351	:	dt	<=	71	;
						10'd352	:	dt	<=	142	;
						10'd353	:	dt	<=	194	;
						10'd354	:	dt	<=	194	;
						10'd355	:	dt	<=	169	;
						10'd356	:	dt	<=	110	;
						10'd357	:	dt	<=	162	;
						10'd358	:	dt	<=	174	;
						10'd359	:	dt	<=	171	;
						10'd360	:	dt	<=	170	;
						10'd361	:	dt	<=	169	;
						10'd362	:	dt	<=	169	;
						10'd363	:	dt	<=	168	;
						10'd364	:	dt	<=	129	;
						10'd365	:	dt	<=	133	;
						10'd366	:	dt	<=	139	;
						10'd367	:	dt	<=	139	;
						10'd368	:	dt	<=	164	;
						10'd369	:	dt	<=	212	;
						10'd370	:	dt	<=	178	;
						10'd371	:	dt	<=	176	;
						10'd372	:	dt	<=	165	;
						10'd373	:	dt	<=	108	;
						10'd374	:	dt	<=	103	;
						10'd375	:	dt	<=	182	;
						10'd376	:	dt	<=	129	;
						10'd377	:	dt	<=	59	;
						10'd378	:	dt	<=	54	;
						10'd379	:	dt	<=	136	;
						10'd380	:	dt	<=	173	;
						10'd381	:	dt	<=	172	;
						10'd382	:	dt	<=	176	;
						10'd383	:	dt	<=	168	;
						10'd384	:	dt	<=	113	;
						10'd385	:	dt	<=	117	;
						10'd386	:	dt	<=	180	;
						10'd387	:	dt	<=	171	;
						10'd388	:	dt	<=	171	;
						10'd389	:	dt	<=	170	;
						10'd390	:	dt	<=	169	;
						10'd391	:	dt	<=	169	;
						10'd392	:	dt	<=	130	;
						10'd393	:	dt	<=	134	;
						10'd394	:	dt	<=	141	;
						10'd395	:	dt	<=	138	;
						10'd396	:	dt	<=	197	;
						10'd397	:	dt	<=	208	;
						10'd398	:	dt	<=	168	;
						10'd399	:	dt	<=	153	;
						10'd400	:	dt	<=	164	;
						10'd401	:	dt	<=	125	;
						10'd402	:	dt	<=	69	;
						10'd403	:	dt	<=	156	;
						10'd404	:	dt	<=	152	;
						10'd405	:	dt	<=	106	;
						10'd406	:	dt	<=	153	;
						10'd407	:	dt	<=	193	;
						10'd408	:	dt	<=	178	;
						10'd409	:	dt	<=	172	;
						10'd410	:	dt	<=	151	;
						10'd411	:	dt	<=	133	;
						10'd412	:	dt	<=	134	;
						10'd413	:	dt	<=	95	;
						10'd414	:	dt	<=	165	;
						10'd415	:	dt	<=	175	;
						10'd416	:	dt	<=	173	;
						10'd417	:	dt	<=	171	;
						10'd418	:	dt	<=	170	;
						10'd419	:	dt	<=	169	;
						10'd420	:	dt	<=	131	;
						10'd421	:	dt	<=	135	;
						10'd422	:	dt	<=	142	;
						10'd423	:	dt	<=	138	;
						10'd424	:	dt	<=	202	;
						10'd425	:	dt	<=	209	;
						10'd426	:	dt	<=	179	;
						10'd427	:	dt	<=	141	;
						10'd428	:	dt	<=	137	;
						10'd429	:	dt	<=	160	;
						10'd430	:	dt	<=	96	;
						10'd431	:	dt	<=	126	;
						10'd432	:	dt	<=	191	;
						10'd433	:	dt	<=	200	;
						10'd434	:	dt	<=	195	;
						10'd435	:	dt	<=	177	;
						10'd436	:	dt	<=	168	;
						10'd437	:	dt	<=	163	;
						10'd438	:	dt	<=	138	;
						10'd439	:	dt	<=	116	;
						10'd440	:	dt	<=	120	;
						10'd441	:	dt	<=	98	;
						10'd442	:	dt	<=	160	;
						10'd443	:	dt	<=	176	;
						10'd444	:	dt	<=	172	;
						10'd445	:	dt	<=	172	;
						10'd446	:	dt	<=	172	;
						10'd447	:	dt	<=	170	;
						10'd448	:	dt	<=	130	;
						10'd449	:	dt	<=	134	;
						10'd450	:	dt	<=	141	;
						10'd451	:	dt	<=	139	;
						10'd452	:	dt	<=	206	;
						10'd453	:	dt	<=	214	;
						10'd454	:	dt	<=	189	;
						10'd455	:	dt	<=	176	;
						10'd456	:	dt	<=	154	;
						10'd457	:	dt	<=	158	;
						10'd458	:	dt	<=	176	;
						10'd459	:	dt	<=	191	;
						10'd460	:	dt	<=	206	;
						10'd461	:	dt	<=	205	;
						10'd462	:	dt	<=	182	;
						10'd463	:	dt	<=	168	;
						10'd464	:	dt	<=	166	;
						10'd465	:	dt	<=	142	;
						10'd466	:	dt	<=	124	;
						10'd467	:	dt	<=	106	;
						10'd468	:	dt	<=	92	;
						10'd469	:	dt	<=	125	;
						10'd470	:	dt	<=	177	;
						10'd471	:	dt	<=	172	;
						10'd472	:	dt	<=	172	;
						10'd473	:	dt	<=	173	;
						10'd474	:	dt	<=	172	;
						10'd475	:	dt	<=	170	;
						10'd476	:	dt	<=	127	;
						10'd477	:	dt	<=	133	;
						10'd478	:	dt	<=	139	;
						10'd479	:	dt	<=	140	;
						10'd480	:	dt	<=	208	;
						10'd481	:	dt	<=	218	;
						10'd482	:	dt	<=	198	;
						10'd483	:	dt	<=	187	;
						10'd484	:	dt	<=	174	;
						10'd485	:	dt	<=	159	;
						10'd486	:	dt	<=	182	;
						10'd487	:	dt	<=	203	;
						10'd488	:	dt	<=	203	;
						10'd489	:	dt	<=	198	;
						10'd490	:	dt	<=	174	;
						10'd491	:	dt	<=	154	;
						10'd492	:	dt	<=	146	;
						10'd493	:	dt	<=	129	;
						10'd494	:	dt	<=	118	;
						10'd495	:	dt	<=	90	;
						10'd496	:	dt	<=	98	;
						10'd497	:	dt	<=	167	;
						10'd498	:	dt	<=	174	;
						10'd499	:	dt	<=	172	;
						10'd500	:	dt	<=	171	;
						10'd501	:	dt	<=	171	;
						10'd502	:	dt	<=	170	;
						10'd503	:	dt	<=	169	;
						10'd504	:	dt	<=	131	;
						10'd505	:	dt	<=	136	;
						10'd506	:	dt	<=	142	;
						10'd507	:	dt	<=	140	;
						10'd508	:	dt	<=	202	;
						10'd509	:	dt	<=	218	;
						10'd510	:	dt	<=	203	;
						10'd511	:	dt	<=	187	;
						10'd512	:	dt	<=	173	;
						10'd513	:	dt	<=	161	;
						10'd514	:	dt	<=	177	;
						10'd515	:	dt	<=	199	;
						10'd516	:	dt	<=	199	;
						10'd517	:	dt	<=	183	;
						10'd518	:	dt	<=	160	;
						10'd519	:	dt	<=	138	;
						10'd520	:	dt	<=	128	;
						10'd521	:	dt	<=	127	;
						10'd522	:	dt	<=	104	;
						10'd523	:	dt	<=	89	;
						10'd524	:	dt	<=	156	;
						10'd525	:	dt	<=	182	;
						10'd526	:	dt	<=	177	;
						10'd527	:	dt	<=	177	;
						10'd528	:	dt	<=	175	;
						10'd529	:	dt	<=	174	;
						10'd530	:	dt	<=	173	;
						10'd531	:	dt	<=	173	;
						10'd532	:	dt	<=	115	;
						10'd533	:	dt	<=	115	;
						10'd534	:	dt	<=	121	;
						10'd535	:	dt	<=	111	;
						10'd536	:	dt	<=	178	;
						10'd537	:	dt	<=	218	;
						10'd538	:	dt	<=	204	;
						10'd539	:	dt	<=	192	;
						10'd540	:	dt	<=	176	;
						10'd541	:	dt	<=	167	;
						10'd542	:	dt	<=	179	;
						10'd543	:	dt	<=	197	;
						10'd544	:	dt	<=	183	;
						10'd545	:	dt	<=	155	;
						10'd546	:	dt	<=	143	;
						10'd547	:	dt	<=	133	;
						10'd548	:	dt	<=	131	;
						10'd549	:	dt	<=	115	;
						10'd550	:	dt	<=	89	;
						10'd551	:	dt	<=	95	;
						10'd552	:	dt	<=	126	;
						10'd553	:	dt	<=	123	;
						10'd554	:	dt	<=	123	;
						10'd555	:	dt	<=	121	;
						10'd556	:	dt	<=	120	;
						10'd557	:	dt	<=	120	;
						10'd558	:	dt	<=	119	;
						10'd559	:	dt	<=	119	;
						10'd560	:	dt	<=	87	;
						10'd561	:	dt	<=	88	;
						10'd562	:	dt	<=	92	;
						10'd563	:	dt	<=	78	;
						10'd564	:	dt	<=	131	;
						10'd565	:	dt	<=	217	;
						10'd566	:	dt	<=	203	;
						10'd567	:	dt	<=	194	;
						10'd568	:	dt	<=	179	;
						10'd569	:	dt	<=	173	;
						10'd570	:	dt	<=	177	;
						10'd571	:	dt	<=	191	;
						10'd572	:	dt	<=	173	;
						10'd573	:	dt	<=	143	;
						10'd574	:	dt	<=	129	;
						10'd575	:	dt	<=	135	;
						10'd576	:	dt	<=	126	;
						10'd577	:	dt	<=	99	;
						10'd578	:	dt	<=	88	;
						10'd579	:	dt	<=	85	;
						10'd580	:	dt	<=	81	;
						10'd581	:	dt	<=	79	;
						10'd582	:	dt	<=	79	;
						10'd583	:	dt	<=	78	;
						10'd584	:	dt	<=	78	;
						10'd585	:	dt	<=	77	;
						10'd586	:	dt	<=	76	;
						10'd587	:	dt	<=	76	;
						10'd588	:	dt	<=	95	;
						10'd589	:	dt	<=	97	;
						10'd590	:	dt	<=	97	;
						10'd591	:	dt	<=	93	;
						10'd592	:	dt	<=	106	;
						10'd593	:	dt	<=	206	;
						10'd594	:	dt	<=	197	;
						10'd595	:	dt	<=	193	;
						10'd596	:	dt	<=	180	;
						10'd597	:	dt	<=	168	;
						10'd598	:	dt	<=	169	;
						10'd599	:	dt	<=	188	;
						10'd600	:	dt	<=	174	;
						10'd601	:	dt	<=	135	;
						10'd602	:	dt	<=	118	;
						10'd603	:	dt	<=	121	;
						10'd604	:	dt	<=	104	;
						10'd605	:	dt	<=	89	;
						10'd606	:	dt	<=	90	;
						10'd607	:	dt	<=	91	;
						10'd608	:	dt	<=	91	;
						10'd609	:	dt	<=	89	;
						10'd610	:	dt	<=	87	;
						10'd611	:	dt	<=	87	;
						10'd612	:	dt	<=	86	;
						10'd613	:	dt	<=	85	;
						10'd614	:	dt	<=	85	;
						10'd615	:	dt	<=	85	;
						10'd616	:	dt	<=	94	;
						10'd617	:	dt	<=	95	;
						10'd618	:	dt	<=	97	;
						10'd619	:	dt	<=	98	;
						10'd620	:	dt	<=	94	;
						10'd621	:	dt	<=	190	;
						10'd622	:	dt	<=	190	;
						10'd623	:	dt	<=	193	;
						10'd624	:	dt	<=	186	;
						10'd625	:	dt	<=	170	;
						10'd626	:	dt	<=	164	;
						10'd627	:	dt	<=	185	;
						10'd628	:	dt	<=	170	;
						10'd629	:	dt	<=	121	;
						10'd630	:	dt	<=	107	;
						10'd631	:	dt	<=	105	;
						10'd632	:	dt	<=	91	;
						10'd633	:	dt	<=	88	;
						10'd634	:	dt	<=	91	;
						10'd635	:	dt	<=	88	;
						10'd636	:	dt	<=	89	;
						10'd637	:	dt	<=	90	;
						10'd638	:	dt	<=	89	;
						10'd639	:	dt	<=	87	;
						10'd640	:	dt	<=	86	;
						10'd641	:	dt	<=	86	;
						10'd642	:	dt	<=	86	;
						10'd643	:	dt	<=	85	;
						10'd644	:	dt	<=	97	;
						10'd645	:	dt	<=	98	;
						10'd646	:	dt	<=	97	;
						10'd647	:	dt	<=	99	;
						10'd648	:	dt	<=	88	;
						10'd649	:	dt	<=	176	;
						10'd650	:	dt	<=	192	;
						10'd651	:	dt	<=	197	;
						10'd652	:	dt	<=	194	;
						10'd653	:	dt	<=	177	;
						10'd654	:	dt	<=	159	;
						10'd655	:	dt	<=	178	;
						10'd656	:	dt	<=	168	;
						10'd657	:	dt	<=	119	;
						10'd658	:	dt	<=	105	;
						10'd659	:	dt	<=	95	;
						10'd660	:	dt	<=	88	;
						10'd661	:	dt	<=	92	;
						10'd662	:	dt	<=	91	;
						10'd663	:	dt	<=	89	;
						10'd664	:	dt	<=	88	;
						10'd665	:	dt	<=	89	;
						10'd666	:	dt	<=	89	;
						10'd667	:	dt	<=	88	;
						10'd668	:	dt	<=	87	;
						10'd669	:	dt	<=	88	;
						10'd670	:	dt	<=	86	;
						10'd671	:	dt	<=	85	;
						10'd672	:	dt	<=	98	;
						10'd673	:	dt	<=	100	;
						10'd674	:	dt	<=	99	;
						10'd675	:	dt	<=	101	;
						10'd676	:	dt	<=	86	;
						10'd677	:	dt	<=	164	;
						10'd678	:	dt	<=	200	;
						10'd679	:	dt	<=	205	;
						10'd680	:	dt	<=	202	;
						10'd681	:	dt	<=	186	;
						10'd682	:	dt	<=	156	;
						10'd683	:	dt	<=	170	;
						10'd684	:	dt	<=	171	;
						10'd685	:	dt	<=	124	;
						10'd686	:	dt	<=	101	;
						10'd687	:	dt	<=	88	;
						10'd688	:	dt	<=	88	;
						10'd689	:	dt	<=	93	;
						10'd690	:	dt	<=	91	;
						10'd691	:	dt	<=	89	;
						10'd692	:	dt	<=	88	;
						10'd693	:	dt	<=	88	;
						10'd694	:	dt	<=	89	;
						10'd695	:	dt	<=	87	;
						10'd696	:	dt	<=	86	;
						10'd697	:	dt	<=	87	;
						10'd698	:	dt	<=	85	;
						10'd699	:	dt	<=	85	;
						10'd700	:	dt	<=	97	;
						10'd701	:	dt	<=	99	;
						10'd702	:	dt	<=	99	;
						10'd703	:	dt	<=	103	;
						10'd704	:	dt	<=	90	;
						10'd705	:	dt	<=	141	;
						10'd706	:	dt	<=	209	;
						10'd707	:	dt	<=	207	;
						10'd708	:	dt	<=	202	;
						10'd709	:	dt	<=	184	;
						10'd710	:	dt	<=	156	;
						10'd711	:	dt	<=	163	;
						10'd712	:	dt	<=	172	;
						10'd713	:	dt	<=	126	;
						10'd714	:	dt	<=	97	;
						10'd715	:	dt	<=	84	;
						10'd716	:	dt	<=	88	;
						10'd717	:	dt	<=	94	;
						10'd718	:	dt	<=	92	;
						10'd719	:	dt	<=	90	;
						10'd720	:	dt	<=	89	;
						10'd721	:	dt	<=	90	;
						10'd722	:	dt	<=	88	;
						10'd723	:	dt	<=	86	;
						10'd724	:	dt	<=	88	;
						10'd725	:	dt	<=	87	;
						10'd726	:	dt	<=	86	;
						10'd727	:	dt	<=	79	;
						10'd728	:	dt	<=	98	;
						10'd729	:	dt	<=	99	;
						10'd730	:	dt	<=	98	;
						10'd731	:	dt	<=	98	;
						10'd732	:	dt	<=	95	;
						10'd733	:	dt	<=	112	;
						10'd734	:	dt	<=	202	;
						10'd735	:	dt	<=	198	;
						10'd736	:	dt	<=	181	;
						10'd737	:	dt	<=	168	;
						10'd738	:	dt	<=	155	;
						10'd739	:	dt	<=	156	;
						10'd740	:	dt	<=	165	;
						10'd741	:	dt	<=	126	;
						10'd742	:	dt	<=	97	;
						10'd743	:	dt	<=	82	;
						10'd744	:	dt	<=	90	;
						10'd745	:	dt	<=	93	;
						10'd746	:	dt	<=	91	;
						10'd747	:	dt	<=	90	;
						10'd748	:	dt	<=	90	;
						10'd749	:	dt	<=	92	;
						10'd750	:	dt	<=	88	;
						10'd751	:	dt	<=	86	;
						10'd752	:	dt	<=	88	;
						10'd753	:	dt	<=	88	;
						10'd754	:	dt	<=	79	;
						10'd755	:	dt	<=	143	;
						10'd756	:	dt	<=	98	;
						10'd757	:	dt	<=	98	;
						10'd758	:	dt	<=	99	;
						10'd759	:	dt	<=	99	;
						10'd760	:	dt	<=	99	;
						10'd761	:	dt	<=	98	;
						10'd762	:	dt	<=	192	;
						10'd763	:	dt	<=	194	;
						10'd764	:	dt	<=	164	;
						10'd765	:	dt	<=	162	;
						10'd766	:	dt	<=	165	;
						10'd767	:	dt	<=	149	;
						10'd768	:	dt	<=	155	;
						10'd769	:	dt	<=	130	;
						10'd770	:	dt	<=	98	;
						10'd771	:	dt	<=	81	;
						10'd772	:	dt	<=	88	;
						10'd773	:	dt	<=	94	;
						10'd774	:	dt	<=	92	;
						10'd775	:	dt	<=	90	;
						10'd776	:	dt	<=	90	;
						10'd777	:	dt	<=	93	;
						10'd778	:	dt	<=	88	;
						10'd779	:	dt	<=	86	;
						10'd780	:	dt	<=	88	;
						10'd781	:	dt	<=	80	;
						10'd782	:	dt	<=	120	;
						10'd783	:	dt	<=	201	;
					endcase
				end
				2'd3	:	begin
					case (cnt)
						10'd0	:	dt	<=	70	;
						10'd1	:	dt	<=	74	;
						10'd2	:	dt	<=	78	;
						10'd3	:	dt	<=	82	;
						10'd4	:	dt	<=	85	;
						10'd5	:	dt	<=	91	;
						10'd6	:	dt	<=	103	;
						10'd7	:	dt	<=	116	;
						10'd8	:	dt	<=	126	;
						10'd9	:	dt	<=	132	;
						10'd10	:	dt	<=	136	;
						10'd11	:	dt	<=	140	;
						10'd12	:	dt	<=	145	;
						10'd13	:	dt	<=	151	;
						10'd14	:	dt	<=	155	;
						10'd15	:	dt	<=	157	;
						10'd16	:	dt	<=	162	;
						10'd17	:	dt	<=	164	;
						10'd18	:	dt	<=	166	;
						10'd19	:	dt	<=	168	;
						10'd20	:	dt	<=	170	;
						10'd21	:	dt	<=	173	;
						10'd22	:	dt	<=	174	;
						10'd23	:	dt	<=	174	;
						10'd24	:	dt	<=	174	;
						10'd25	:	dt	<=	175	;
						10'd26	:	dt	<=	176	;
						10'd27	:	dt	<=	175	;
						10'd28	:	dt	<=	72	;
						10'd29	:	dt	<=	75	;
						10'd30	:	dt	<=	77	;
						10'd31	:	dt	<=	83	;
						10'd32	:	dt	<=	86	;
						10'd33	:	dt	<=	91	;
						10'd34	:	dt	<=	104	;
						10'd35	:	dt	<=	117	;
						10'd36	:	dt	<=	126	;
						10'd37	:	dt	<=	134	;
						10'd38	:	dt	<=	138	;
						10'd39	:	dt	<=	140	;
						10'd40	:	dt	<=	146	;
						10'd41	:	dt	<=	151	;
						10'd42	:	dt	<=	155	;
						10'd43	:	dt	<=	159	;
						10'd44	:	dt	<=	163	;
						10'd45	:	dt	<=	166	;
						10'd46	:	dt	<=	168	;
						10'd47	:	dt	<=	171	;
						10'd48	:	dt	<=	173	;
						10'd49	:	dt	<=	173	;
						10'd50	:	dt	<=	176	;
						10'd51	:	dt	<=	176	;
						10'd52	:	dt	<=	175	;
						10'd53	:	dt	<=	178	;
						10'd54	:	dt	<=	180	;
						10'd55	:	dt	<=	179	;
						10'd56	:	dt	<=	72	;
						10'd57	:	dt	<=	74	;
						10'd58	:	dt	<=	77	;
						10'd59	:	dt	<=	83	;
						10'd60	:	dt	<=	89	;
						10'd61	:	dt	<=	94	;
						10'd62	:	dt	<=	108	;
						10'd63	:	dt	<=	119	;
						10'd64	:	dt	<=	128	;
						10'd65	:	dt	<=	136	;
						10'd66	:	dt	<=	141	;
						10'd67	:	dt	<=	142	;
						10'd68	:	dt	<=	148	;
						10'd69	:	dt	<=	155	;
						10'd70	:	dt	<=	158	;
						10'd71	:	dt	<=	163	;
						10'd72	:	dt	<=	166	;
						10'd73	:	dt	<=	169	;
						10'd74	:	dt	<=	170	;
						10'd75	:	dt	<=	172	;
						10'd76	:	dt	<=	174	;
						10'd77	:	dt	<=	176	;
						10'd78	:	dt	<=	177	;
						10'd79	:	dt	<=	179	;
						10'd80	:	dt	<=	180	;
						10'd81	:	dt	<=	179	;
						10'd82	:	dt	<=	180	;
						10'd83	:	dt	<=	180	;
						10'd84	:	dt	<=	73	;
						10'd85	:	dt	<=	75	;
						10'd86	:	dt	<=	78	;
						10'd87	:	dt	<=	85	;
						10'd88	:	dt	<=	82	;
						10'd89	:	dt	<=	89	;
						10'd90	:	dt	<=	106	;
						10'd91	:	dt	<=	119	;
						10'd92	:	dt	<=	128	;
						10'd93	:	dt	<=	136	;
						10'd94	:	dt	<=	141	;
						10'd95	:	dt	<=	144	;
						10'd96	:	dt	<=	149	;
						10'd97	:	dt	<=	156	;
						10'd98	:	dt	<=	159	;
						10'd99	:	dt	<=	164	;
						10'd100	:	dt	<=	168	;
						10'd101	:	dt	<=	170	;
						10'd102	:	dt	<=	172	;
						10'd103	:	dt	<=	175	;
						10'd104	:	dt	<=	177	;
						10'd105	:	dt	<=	179	;
						10'd106	:	dt	<=	179	;
						10'd107	:	dt	<=	181	;
						10'd108	:	dt	<=	183	;
						10'd109	:	dt	<=	181	;
						10'd110	:	dt	<=	181	;
						10'd111	:	dt	<=	182	;
						10'd112	:	dt	<=	73	;
						10'd113	:	dt	<=	75	;
						10'd114	:	dt	<=	79	;
						10'd115	:	dt	<=	81	;
						10'd116	:	dt	<=	118	;
						10'd117	:	dt	<=	127	;
						10'd118	:	dt	<=	126	;
						10'd119	:	dt	<=	126	;
						10'd120	:	dt	<=	135	;
						10'd121	:	dt	<=	143	;
						10'd122	:	dt	<=	142	;
						10'd123	:	dt	<=	146	;
						10'd124	:	dt	<=	151	;
						10'd125	:	dt	<=	158	;
						10'd126	:	dt	<=	164	;
						10'd127	:	dt	<=	166	;
						10'd128	:	dt	<=	167	;
						10'd129	:	dt	<=	170	;
						10'd130	:	dt	<=	174	;
						10'd131	:	dt	<=	177	;
						10'd132	:	dt	<=	179	;
						10'd133	:	dt	<=	181	;
						10'd134	:	dt	<=	181	;
						10'd135	:	dt	<=	183	;
						10'd136	:	dt	<=	186	;
						10'd137	:	dt	<=	185	;
						10'd138	:	dt	<=	185	;
						10'd139	:	dt	<=	186	;
						10'd140	:	dt	<=	72	;
						10'd141	:	dt	<=	79	;
						10'd142	:	dt	<=	69	;
						10'd143	:	dt	<=	127	;
						10'd144	:	dt	<=	208	;
						10'd145	:	dt	<=	148	;
						10'd146	:	dt	<=	139	;
						10'd147	:	dt	<=	133	;
						10'd148	:	dt	<=	151	;
						10'd149	:	dt	<=	162	;
						10'd150	:	dt	<=	144	;
						10'd151	:	dt	<=	138	;
						10'd152	:	dt	<=	140	;
						10'd153	:	dt	<=	151	;
						10'd154	:	dt	<=	153	;
						10'd155	:	dt	<=	165	;
						10'd156	:	dt	<=	175	;
						10'd157	:	dt	<=	176	;
						10'd158	:	dt	<=	178	;
						10'd159	:	dt	<=	178	;
						10'd160	:	dt	<=	180	;
						10'd161	:	dt	<=	183	;
						10'd162	:	dt	<=	185	;
						10'd163	:	dt	<=	187	;
						10'd164	:	dt	<=	187	;
						10'd165	:	dt	<=	187	;
						10'd166	:	dt	<=	187	;
						10'd167	:	dt	<=	187	;
						10'd168	:	dt	<=	74	;
						10'd169	:	dt	<=	80	;
						10'd170	:	dt	<=	69	;
						10'd171	:	dt	<=	127	;
						10'd172	:	dt	<=	173	;
						10'd173	:	dt	<=	104	;
						10'd174	:	dt	<=	104	;
						10'd175	:	dt	<=	102	;
						10'd176	:	dt	<=	144	;
						10'd177	:	dt	<=	142	;
						10'd178	:	dt	<=	120	;
						10'd179	:	dt	<=	121	;
						10'd180	:	dt	<=	163	;
						10'd181	:	dt	<=	164	;
						10'd182	:	dt	<=	136	;
						10'd183	:	dt	<=	124	;
						10'd184	:	dt	<=	136	;
						10'd185	:	dt	<=	161	;
						10'd186	:	dt	<=	172	;
						10'd187	:	dt	<=	184	;
						10'd188	:	dt	<=	187	;
						10'd189	:	dt	<=	183	;
						10'd190	:	dt	<=	186	;
						10'd191	:	dt	<=	189	;
						10'd192	:	dt	<=	189	;
						10'd193	:	dt	<=	189	;
						10'd194	:	dt	<=	189	;
						10'd195	:	dt	<=	189	;
						10'd196	:	dt	<=	75	;
						10'd197	:	dt	<=	76	;
						10'd198	:	dt	<=	79	;
						10'd199	:	dt	<=	83	;
						10'd200	:	dt	<=	99	;
						10'd201	:	dt	<=	90	;
						10'd202	:	dt	<=	93	;
						10'd203	:	dt	<=	89	;
						10'd204	:	dt	<=	125	;
						10'd205	:	dt	<=	116	;
						10'd206	:	dt	<=	96	;
						10'd207	:	dt	<=	109	;
						10'd208	:	dt	<=	168	;
						10'd209	:	dt	<=	168	;
						10'd210	:	dt	<=	145	;
						10'd211	:	dt	<=	104	;
						10'd212	:	dt	<=	123	;
						10'd213	:	dt	<=	133	;
						10'd214	:	dt	<=	142	;
						10'd215	:	dt	<=	138	;
						10'd216	:	dt	<=	165	;
						10'd217	:	dt	<=	194	;
						10'd218	:	dt	<=	186	;
						10'd219	:	dt	<=	190	;
						10'd220	:	dt	<=	191	;
						10'd221	:	dt	<=	190	;
						10'd222	:	dt	<=	191	;
						10'd223	:	dt	<=	190	;
						10'd224	:	dt	<=	75	;
						10'd225	:	dt	<=	77	;
						10'd226	:	dt	<=	81	;
						10'd227	:	dt	<=	85	;
						10'd228	:	dt	<=	86	;
						10'd229	:	dt	<=	98	;
						10'd230	:	dt	<=	110	;
						10'd231	:	dt	<=	118	;
						10'd232	:	dt	<=	125	;
						10'd233	:	dt	<=	121	;
						10'd234	:	dt	<=	111	;
						10'd235	:	dt	<=	114	;
						10'd236	:	dt	<=	155	;
						10'd237	:	dt	<=	160	;
						10'd238	:	dt	<=	118	;
						10'd239	:	dt	<=	109	;
						10'd240	:	dt	<=	170	;
						10'd241	:	dt	<=	151	;
						10'd242	:	dt	<=	149	;
						10'd243	:	dt	<=	136	;
						10'd244	:	dt	<=	98	;
						10'd245	:	dt	<=	155	;
						10'd246	:	dt	<=	200	;
						10'd247	:	dt	<=	189	;
						10'd248	:	dt	<=	194	;
						10'd249	:	dt	<=	192	;
						10'd250	:	dt	<=	193	;
						10'd251	:	dt	<=	192	;
						10'd252	:	dt	<=	75	;
						10'd253	:	dt	<=	78	;
						10'd254	:	dt	<=	81	;
						10'd255	:	dt	<=	85	;
						10'd256	:	dt	<=	89	;
						10'd257	:	dt	<=	99	;
						10'd258	:	dt	<=	115	;
						10'd259	:	dt	<=	129	;
						10'd260	:	dt	<=	140	;
						10'd261	:	dt	<=	148	;
						10'd262	:	dt	<=	148	;
						10'd263	:	dt	<=	148	;
						10'd264	:	dt	<=	140	;
						10'd265	:	dt	<=	114	;
						10'd266	:	dt	<=	91	;
						10'd267	:	dt	<=	194	;
						10'd268	:	dt	<=	164	;
						10'd269	:	dt	<=	164	;
						10'd270	:	dt	<=	126	;
						10'd271	:	dt	<=	165	;
						10'd272	:	dt	<=	139	;
						10'd273	:	dt	<=	82	;
						10'd274	:	dt	<=	169	;
						10'd275	:	dt	<=	200	;
						10'd276	:	dt	<=	193	;
						10'd277	:	dt	<=	195	;
						10'd278	:	dt	<=	196	;
						10'd279	:	dt	<=	195	;
						10'd280	:	dt	<=	77	;
						10'd281	:	dt	<=	77	;
						10'd282	:	dt	<=	81	;
						10'd283	:	dt	<=	85	;
						10'd284	:	dt	<=	88	;
						10'd285	:	dt	<=	100	;
						10'd286	:	dt	<=	115	;
						10'd287	:	dt	<=	128	;
						10'd288	:	dt	<=	139	;
						10'd289	:	dt	<=	144	;
						10'd290	:	dt	<=	155	;
						10'd291	:	dt	<=	190	;
						10'd292	:	dt	<=	127	;
						10'd293	:	dt	<=	92	;
						10'd294	:	dt	<=	100	;
						10'd295	:	dt	<=	167	;
						10'd296	:	dt	<=	158	;
						10'd297	:	dt	<=	123	;
						10'd298	:	dt	<=	122	;
						10'd299	:	dt	<=	165	;
						10'd300	:	dt	<=	144	;
						10'd301	:	dt	<=	125	;
						10'd302	:	dt	<=	76	;
						10'd303	:	dt	<=	187	;
						10'd304	:	dt	<=	198	;
						10'd305	:	dt	<=	195	;
						10'd306	:	dt	<=	196	;
						10'd307	:	dt	<=	196	;
						10'd308	:	dt	<=	75	;
						10'd309	:	dt	<=	77	;
						10'd310	:	dt	<=	80	;
						10'd311	:	dt	<=	85	;
						10'd312	:	dt	<=	88	;
						10'd313	:	dt	<=	101	;
						10'd314	:	dt	<=	116	;
						10'd315	:	dt	<=	129	;
						10'd316	:	dt	<=	141	;
						10'd317	:	dt	<=	143	;
						10'd318	:	dt	<=	176	;
						10'd319	:	dt	<=	201	;
						10'd320	:	dt	<=	159	;
						10'd321	:	dt	<=	91	;
						10'd322	:	dt	<=	66	;
						10'd323	:	dt	<=	68	;
						10'd324	:	dt	<=	111	;
						10'd325	:	dt	<=	91	;
						10'd326	:	dt	<=	148	;
						10'd327	:	dt	<=	129	;
						10'd328	:	dt	<=	135	;
						10'd329	:	dt	<=	146	;
						10'd330	:	dt	<=	79	;
						10'd331	:	dt	<=	98	;
						10'd332	:	dt	<=	208	;
						10'd333	:	dt	<=	196	;
						10'd334	:	dt	<=	198	;
						10'd335	:	dt	<=	198	;
						10'd336	:	dt	<=	76	;
						10'd337	:	dt	<=	78	;
						10'd338	:	dt	<=	81	;
						10'd339	:	dt	<=	84	;
						10'd340	:	dt	<=	88	;
						10'd341	:	dt	<=	101	;
						10'd342	:	dt	<=	118	;
						10'd343	:	dt	<=	130	;
						10'd344	:	dt	<=	141	;
						10'd345	:	dt	<=	145	;
						10'd346	:	dt	<=	164	;
						10'd347	:	dt	<=	205	;
						10'd348	:	dt	<=	189	;
						10'd349	:	dt	<=	138	;
						10'd350	:	dt	<=	114	;
						10'd351	:	dt	<=	92	;
						10'd352	:	dt	<=	77	;
						10'd353	:	dt	<=	95	;
						10'd354	:	dt	<=	167	;
						10'd355	:	dt	<=	124	;
						10'd356	:	dt	<=	135	;
						10'd357	:	dt	<=	106	;
						10'd358	:	dt	<=	101	;
						10'd359	:	dt	<=	54	;
						10'd360	:	dt	<=	147	;
						10'd361	:	dt	<=	214	;
						10'd362	:	dt	<=	197	;
						10'd363	:	dt	<=	200	;
						10'd364	:	dt	<=	75	;
						10'd365	:	dt	<=	78	;
						10'd366	:	dt	<=	80	;
						10'd367	:	dt	<=	84	;
						10'd368	:	dt	<=	89	;
						10'd369	:	dt	<=	102	;
						10'd370	:	dt	<=	119	;
						10'd371	:	dt	<=	130	;
						10'd372	:	dt	<=	141	;
						10'd373	:	dt	<=	147	;
						10'd374	:	dt	<=	178	;
						10'd375	:	dt	<=	175	;
						10'd376	:	dt	<=	183	;
						10'd377	:	dt	<=	166	;
						10'd378	:	dt	<=	183	;
						10'd379	:	dt	<=	158	;
						10'd380	:	dt	<=	96	;
						10'd381	:	dt	<=	94	;
						10'd382	:	dt	<=	93	;
						10'd383	:	dt	<=	102	;
						10'd384	:	dt	<=	101	;
						10'd385	:	dt	<=	71	;
						10'd386	:	dt	<=	60	;
						10'd387	:	dt	<=	64	;
						10'd388	:	dt	<=	59	;
						10'd389	:	dt	<=	186	;
						10'd390	:	dt	<=	207	;
						10'd391	:	dt	<=	200	;
						10'd392	:	dt	<=	76	;
						10'd393	:	dt	<=	78	;
						10'd394	:	dt	<=	80	;
						10'd395	:	dt	<=	85	;
						10'd396	:	dt	<=	89	;
						10'd397	:	dt	<=	102	;
						10'd398	:	dt	<=	117	;
						10'd399	:	dt	<=	132	;
						10'd400	:	dt	<=	138	;
						10'd401	:	dt	<=	166	;
						10'd402	:	dt	<=	196	;
						10'd403	:	dt	<=	158	;
						10'd404	:	dt	<=	156	;
						10'd405	:	dt	<=	140	;
						10'd406	:	dt	<=	178	;
						10'd407	:	dt	<=	150	;
						10'd408	:	dt	<=	77	;
						10'd409	:	dt	<=	78	;
						10'd410	:	dt	<=	82	;
						10'd411	:	dt	<=	75	;
						10'd412	:	dt	<=	87	;
						10'd413	:	dt	<=	68	;
						10'd414	:	dt	<=	47	;
						10'd415	:	dt	<=	57	;
						10'd416	:	dt	<=	44	;
						10'd417	:	dt	<=	75	;
						10'd418	:	dt	<=	202	;
						10'd419	:	dt	<=	204	;
						10'd420	:	dt	<=	77	;
						10'd421	:	dt	<=	78	;
						10'd422	:	dt	<=	81	;
						10'd423	:	dt	<=	85	;
						10'd424	:	dt	<=	89	;
						10'd425	:	dt	<=	103	;
						10'd426	:	dt	<=	119	;
						10'd427	:	dt	<=	132	;
						10'd428	:	dt	<=	141	;
						10'd429	:	dt	<=	163	;
						10'd430	:	dt	<=	160	;
						10'd431	:	dt	<=	118	;
						10'd432	:	dt	<=	123	;
						10'd433	:	dt	<=	130	;
						10'd434	:	dt	<=	157	;
						10'd435	:	dt	<=	111	;
						10'd436	:	dt	<=	72	;
						10'd437	:	dt	<=	79	;
						10'd438	:	dt	<=	77	;
						10'd439	:	dt	<=	80	;
						10'd440	:	dt	<=	90	;
						10'd441	:	dt	<=	79	;
						10'd442	:	dt	<=	56	;
						10'd443	:	dt	<=	55	;
						10'd444	:	dt	<=	55	;
						10'd445	:	dt	<=	33	;
						10'd446	:	dt	<=	116	;
						10'd447	:	dt	<=	217	;
						10'd448	:	dt	<=	77	;
						10'd449	:	dt	<=	78	;
						10'd450	:	dt	<=	80	;
						10'd451	:	dt	<=	85	;
						10'd452	:	dt	<=	89	;
						10'd453	:	dt	<=	104	;
						10'd454	:	dt	<=	119	;
						10'd455	:	dt	<=	131	;
						10'd456	:	dt	<=	143	;
						10'd457	:	dt	<=	155	;
						10'd458	:	dt	<=	170	;
						10'd459	:	dt	<=	128	;
						10'd460	:	dt	<=	125	;
						10'd461	:	dt	<=	94	;
						10'd462	:	dt	<=	79	;
						10'd463	:	dt	<=	69	;
						10'd464	:	dt	<=	60	;
						10'd465	:	dt	<=	67	;
						10'd466	:	dt	<=	68	;
						10'd467	:	dt	<=	70	;
						10'd468	:	dt	<=	76	;
						10'd469	:	dt	<=	71	;
						10'd470	:	dt	<=	71	;
						10'd471	:	dt	<=	67	;
						10'd472	:	dt	<=	54	;
						10'd473	:	dt	<=	51	;
						10'd474	:	dt	<=	50	;
						10'd475	:	dt	<=	190	;
						10'd476	:	dt	<=	77	;
						10'd477	:	dt	<=	78	;
						10'd478	:	dt	<=	80	;
						10'd479	:	dt	<=	85	;
						10'd480	:	dt	<=	89	;
						10'd481	:	dt	<=	105	;
						10'd482	:	dt	<=	121	;
						10'd483	:	dt	<=	133	;
						10'd484	:	dt	<=	141	;
						10'd485	:	dt	<=	162	;
						10'd486	:	dt	<=	187	;
						10'd487	:	dt	<=	186	;
						10'd488	:	dt	<=	156	;
						10'd489	:	dt	<=	106	;
						10'd490	:	dt	<=	82	;
						10'd491	:	dt	<=	106	;
						10'd492	:	dt	<=	92	;
						10'd493	:	dt	<=	42	;
						10'd494	:	dt	<=	72	;
						10'd495	:	dt	<=	85	;
						10'd496	:	dt	<=	82	;
						10'd497	:	dt	<=	77	;
						10'd498	:	dt	<=	85	;
						10'd499	:	dt	<=	82	;
						10'd500	:	dt	<=	62	;
						10'd501	:	dt	<=	55	;
						10'd502	:	dt	<=	41	;
						10'd503	:	dt	<=	116	;
						10'd504	:	dt	<=	76	;
						10'd505	:	dt	<=	78	;
						10'd506	:	dt	<=	81	;
						10'd507	:	dt	<=	84	;
						10'd508	:	dt	<=	89	;
						10'd509	:	dt	<=	105	;
						10'd510	:	dt	<=	120	;
						10'd511	:	dt	<=	133	;
						10'd512	:	dt	<=	145	;
						10'd513	:	dt	<=	153	;
						10'd514	:	dt	<=	165	;
						10'd515	:	dt	<=	185	;
						10'd516	:	dt	<=	165	;
						10'd517	:	dt	<=	128	;
						10'd518	:	dt	<=	120	;
						10'd519	:	dt	<=	112	;
						10'd520	:	dt	<=	118	;
						10'd521	:	dt	<=	49	;
						10'd522	:	dt	<=	76	;
						10'd523	:	dt	<=	108	;
						10'd524	:	dt	<=	100	;
						10'd525	:	dt	<=	101	;
						10'd526	:	dt	<=	107	;
						10'd527	:	dt	<=	96	;
						10'd528	:	dt	<=	65	;
						10'd529	:	dt	<=	48	;
						10'd530	:	dt	<=	54	;
						10'd531	:	dt	<=	50	;
						10'd532	:	dt	<=	77	;
						10'd533	:	dt	<=	78	;
						10'd534	:	dt	<=	80	;
						10'd535	:	dt	<=	84	;
						10'd536	:	dt	<=	89	;
						10'd537	:	dt	<=	106	;
						10'd538	:	dt	<=	120	;
						10'd539	:	dt	<=	134	;
						10'd540	:	dt	<=	146	;
						10'd541	:	dt	<=	152	;
						10'd542	:	dt	<=	159	;
						10'd543	:	dt	<=	158	;
						10'd544	:	dt	<=	140	;
						10'd545	:	dt	<=	112	;
						10'd546	:	dt	<=	73	;
						10'd547	:	dt	<=	68	;
						10'd548	:	dt	<=	109	;
						10'd549	:	dt	<=	135	;
						10'd550	:	dt	<=	70	;
						10'd551	:	dt	<=	107	;
						10'd552	:	dt	<=	122	;
						10'd553	:	dt	<=	119	;
						10'd554	:	dt	<=	109	;
						10'd555	:	dt	<=	88	;
						10'd556	:	dt	<=	55	;
						10'd557	:	dt	<=	52	;
						10'd558	:	dt	<=	58	;
						10'd559	:	dt	<=	54	;
						10'd560	:	dt	<=	77	;
						10'd561	:	dt	<=	76	;
						10'd562	:	dt	<=	79	;
						10'd563	:	dt	<=	83	;
						10'd564	:	dt	<=	89	;
						10'd565	:	dt	<=	105	;
						10'd566	:	dt	<=	121	;
						10'd567	:	dt	<=	136	;
						10'd568	:	dt	<=	146	;
						10'd569	:	dt	<=	153	;
						10'd570	:	dt	<=	154	;
						10'd571	:	dt	<=	157	;
						10'd572	:	dt	<=	136	;
						10'd573	:	dt	<=	107	;
						10'd574	:	dt	<=	72	;
						10'd575	:	dt	<=	52	;
						10'd576	:	dt	<=	89	;
						10'd577	:	dt	<=	125	;
						10'd578	:	dt	<=	80	;
						10'd579	:	dt	<=	80	;
						10'd580	:	dt	<=	131	;
						10'd581	:	dt	<=	127	;
						10'd582	:	dt	<=	98	;
						10'd583	:	dt	<=	71	;
						10'd584	:	dt	<=	53	;
						10'd585	:	dt	<=	58	;
						10'd586	:	dt	<=	61	;
						10'd587	:	dt	<=	59	;
						10'd588	:	dt	<=	77	;
						10'd589	:	dt	<=	76	;
						10'd590	:	dt	<=	79	;
						10'd591	:	dt	<=	82	;
						10'd592	:	dt	<=	89	;
						10'd593	:	dt	<=	105	;
						10'd594	:	dt	<=	122	;
						10'd595	:	dt	<=	136	;
						10'd596	:	dt	<=	146	;
						10'd597	:	dt	<=	152	;
						10'd598	:	dt	<=	154	;
						10'd599	:	dt	<=	162	;
						10'd600	:	dt	<=	172	;
						10'd601	:	dt	<=	178	;
						10'd602	:	dt	<=	180	;
						10'd603	:	dt	<=	157	;
						10'd604	:	dt	<=	118	;
						10'd605	:	dt	<=	147	;
						10'd606	:	dt	<=	148	;
						10'd607	:	dt	<=	113	;
						10'd608	:	dt	<=	109	;
						10'd609	:	dt	<=	105	;
						10'd610	:	dt	<=	77	;
						10'd611	:	dt	<=	65	;
						10'd612	:	dt	<=	61	;
						10'd613	:	dt	<=	65	;
						10'd614	:	dt	<=	65	;
						10'd615	:	dt	<=	59	;
						10'd616	:	dt	<=	73	;
						10'd617	:	dt	<=	74	;
						10'd618	:	dt	<=	78	;
						10'd619	:	dt	<=	79	;
						10'd620	:	dt	<=	87	;
						10'd621	:	dt	<=	104	;
						10'd622	:	dt	<=	120	;
						10'd623	:	dt	<=	134	;
						10'd624	:	dt	<=	146	;
						10'd625	:	dt	<=	152	;
						10'd626	:	dt	<=	154	;
						10'd627	:	dt	<=	159	;
						10'd628	:	dt	<=	167	;
						10'd629	:	dt	<=	171	;
						10'd630	:	dt	<=	183	;
						10'd631	:	dt	<=	180	;
						10'd632	:	dt	<=	87	;
						10'd633	:	dt	<=	110	;
						10'd634	:	dt	<=	128	;
						10'd635	:	dt	<=	141	;
						10'd636	:	dt	<=	96	;
						10'd637	:	dt	<=	98	;
						10'd638	:	dt	<=	84	;
						10'd639	:	dt	<=	56	;
						10'd640	:	dt	<=	39	;
						10'd641	:	dt	<=	38	;
						10'd642	:	dt	<=	38	;
						10'd643	:	dt	<=	42	;
						10'd644	:	dt	<=	71	;
						10'd645	:	dt	<=	73	;
						10'd646	:	dt	<=	77	;
						10'd647	:	dt	<=	77	;
						10'd648	:	dt	<=	86	;
						10'd649	:	dt	<=	105	;
						10'd650	:	dt	<=	121	;
						10'd651	:	dt	<=	134	;
						10'd652	:	dt	<=	146	;
						10'd653	:	dt	<=	151	;
						10'd654	:	dt	<=	153	;
						10'd655	:	dt	<=	160	;
						10'd656	:	dt	<=	168	;
						10'd657	:	dt	<=	173	;
						10'd658	:	dt	<=	187	;
						10'd659	:	dt	<=	152	;
						10'd660	:	dt	<=	61	;
						10'd661	:	dt	<=	57	;
						10'd662	:	dt	<=	33	;
						10'd663	:	dt	<=	38	;
						10'd664	:	dt	<=	48	;
						10'd665	:	dt	<=	51	;
						10'd666	:	dt	<=	37	;
						10'd667	:	dt	<=	20	;
						10'd668	:	dt	<=	10	;
						10'd669	:	dt	<=	7	;
						10'd670	:	dt	<=	3	;
						10'd671	:	dt	<=	0	;
						10'd672	:	dt	<=	72	;
						10'd673	:	dt	<=	72	;
						10'd674	:	dt	<=	76	;
						10'd675	:	dt	<=	77	;
						10'd676	:	dt	<=	84	;
						10'd677	:	dt	<=	103	;
						10'd678	:	dt	<=	119	;
						10'd679	:	dt	<=	134	;
						10'd680	:	dt	<=	146	;
						10'd681	:	dt	<=	151	;
						10'd682	:	dt	<=	154	;
						10'd683	:	dt	<=	161	;
						10'd684	:	dt	<=	168	;
						10'd685	:	dt	<=	173	;
						10'd686	:	dt	<=	191	;
						10'd687	:	dt	<=	125	;
						10'd688	:	dt	<=	62	;
						10'd689	:	dt	<=	67	;
						10'd690	:	dt	<=	63	;
						10'd691	:	dt	<=	9	;
						10'd692	:	dt	<=	14	;
						10'd693	:	dt	<=	28	;
						10'd694	:	dt	<=	20	;
						10'd695	:	dt	<=	13	;
						10'd696	:	dt	<=	12	;
						10'd697	:	dt	<=	8	;
						10'd698	:	dt	<=	1	;
						10'd699	:	dt	<=	0	;
						10'd700	:	dt	<=	70	;
						10'd701	:	dt	<=	71	;
						10'd702	:	dt	<=	74	;
						10'd703	:	dt	<=	77	;
						10'd704	:	dt	<=	83	;
						10'd705	:	dt	<=	101	;
						10'd706	:	dt	<=	120	;
						10'd707	:	dt	<=	134	;
						10'd708	:	dt	<=	145	;
						10'd709	:	dt	<=	153	;
						10'd710	:	dt	<=	155	;
						10'd711	:	dt	<=	162	;
						10'd712	:	dt	<=	169	;
						10'd713	:	dt	<=	176	;
						10'd714	:	dt	<=	186	;
						10'd715	:	dt	<=	100	;
						10'd716	:	dt	<=	60	;
						10'd717	:	dt	<=	57	;
						10'd718	:	dt	<=	58	;
						10'd719	:	dt	<=	49	;
						10'd720	:	dt	<=	0	;
						10'd721	:	dt	<=	16	;
						10'd722	:	dt	<=	22	;
						10'd723	:	dt	<=	15	;
						10'd724	:	dt	<=	12	;
						10'd725	:	dt	<=	8	;
						10'd726	:	dt	<=	1	;
						10'd727	:	dt	<=	0	;
						10'd728	:	dt	<=	68	;
						10'd729	:	dt	<=	68	;
						10'd730	:	dt	<=	72	;
						10'd731	:	dt	<=	74	;
						10'd732	:	dt	<=	82	;
						10'd733	:	dt	<=	101	;
						10'd734	:	dt	<=	118	;
						10'd735	:	dt	<=	133	;
						10'd736	:	dt	<=	145	;
						10'd737	:	dt	<=	152	;
						10'd738	:	dt	<=	155	;
						10'd739	:	dt	<=	161	;
						10'd740	:	dt	<=	168	;
						10'd741	:	dt	<=	180	;
						10'd742	:	dt	<=	167	;
						10'd743	:	dt	<=	68	;
						10'd744	:	dt	<=	59	;
						10'd745	:	dt	<=	56	;
						10'd746	:	dt	<=	50	;
						10'd747	:	dt	<=	59	;
						10'd748	:	dt	<=	0	;
						10'd749	:	dt	<=	0	;
						10'd750	:	dt	<=	14	;
						10'd751	:	dt	<=	10	;
						10'd752	:	dt	<=	1	;
						10'd753	:	dt	<=	0	;
						10'd754	:	dt	<=	0	;
						10'd755	:	dt	<=	0	;
						10'd756	:	dt	<=	64	;
						10'd757	:	dt	<=	65	;
						10'd758	:	dt	<=	70	;
						10'd759	:	dt	<=	72	;
						10'd760	:	dt	<=	81	;
						10'd761	:	dt	<=	99	;
						10'd762	:	dt	<=	115	;
						10'd763	:	dt	<=	130	;
						10'd764	:	dt	<=	142	;
						10'd765	:	dt	<=	150	;
						10'd766	:	dt	<=	152	;
						10'd767	:	dt	<=	160	;
						10'd768	:	dt	<=	166	;
						10'd769	:	dt	<=	184	;
						10'd770	:	dt	<=	132	;
						10'd771	:	dt	<=	58	;
						10'd772	:	dt	<=	64	;
						10'd773	:	dt	<=	52	;
						10'd774	:	dt	<=	49	;
						10'd775	:	dt	<=	62	;
						10'd776	:	dt	<=	0	;
						10'd777	:	dt	<=	0	;
						10'd778	:	dt	<=	0	;
						10'd779	:	dt	<=	3	;
						10'd780	:	dt	<=	0	;
						10'd781	:	dt	<=	1	;
						10'd782	:	dt	<=	4	;
						10'd783	:	dt	<=	0	;
					endcase
				end
			endcase
		end
	end

	assign	q_data = dt;
	
endmodule
