`include "global.sv"
`include "timescale.sv"

module src_rom(
	input			clk,
	input			rstn,
	input	[11:0]		aa,
	input			cena,
	output reg		[`WD:0]	qa
	);
	logic [0:28*28-1][`WD:0] mem = {			   
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd1,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,
16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0,	16'd0
		   };
		
	always @(posedge clk, negedge rstn)
		if (rstn == 0)	qa <= 0;
		else if (!cena)		qa <= mem[aa];
endmodule