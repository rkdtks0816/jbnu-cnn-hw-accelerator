`include "global.sv"
`include "timescale.sv"
module bias_fc1_rom(
	input			clk,
	input							rstn,
	input	[`W_OUTPUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_FC1 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC1-1][0:`OUTPUT_NUM_FC1-1][`WD_BIAS:0] weight	 = {
-34'd43163716,  34'd170595872,  -34'd296727040,  34'd9611279,  34'd323266912,  -34'd89451704,  34'd605244352,  -34'd410449632,  -34'd10538601,  34'd22564342,  -34'd424003744,  -34'd121739336,  34'd199549760,  34'd442508736,  -34'd566966656,  -34'd17477802,  
-34'd92106680,  34'd457087200,  34'd753293504,  -34'd281958976,  -34'd179784064,  -34'd71860232,  -34'd75914824,  34'd10182526,  -34'd43681848,  -34'd247113520,  -34'd3423327,  34'd306645376,  34'd635585984,  -34'd127214352,  -34'd77502560,  34'd217642112,  
-34'd70771200,  -34'd205134912,  34'd151931888,  -34'd57247372,  34'd135403136,  34'd404339648,  -34'd4743681,  -34'd308377728,  34'd29545812,  -34'd426148864,  -34'd3681535,  -34'd75140896,  -34'd182082112,  -34'd22870048,  34'd158906624,  -34'd208246784,  
34'd582799168,  -34'd302631456,  -34'd197160960,  34'd387801696,  -34'd333398976,  -34'd7022893,  34'd58144684,  -34'd100847408,  34'd401725728,  -34'd194834976,  34'd36175244,  34'd92399064,  34'd273416992,  34'd158028400,  -34'd53797476,  -34'd32233150
	};
	
	always @(posedge clk) begin
		if (rstn == 0) begin
			qa <= 0;
		end
		else if (!cena) begin
			qa <= weight[aa];	
		end
	end
endmodule


