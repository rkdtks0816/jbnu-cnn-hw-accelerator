`include "global.sv"
`include "timescale.sv"

module sign_mnist(
	input							clk,
	input							rstn,
	input							en,
	input							key_1,
	input							iready,
	input				[5:0]		io,
	
	output	reg				ready,
	output			[`WD:0]	q_data,
	output	reg				push
	);
	reg	[`WD:0]		dt;
	
	reg	[1:0]		din;
	reg	[1:0]		rin;
	reg	[1:0]		rpush;
	reg	[4:0]		count;
	
	reg	[10:0]		cnt;
	reg					cnt_en;
	wire			cnt_max = cnt == 10'd783;
	wire			end_cnt_en = cnt_max;
	

	always @(posedge clk, negedge rstn) begin
		if(rstn == 0) begin
			din	<=	2'd0;
			push	<=	1'b0;
		end
		else begin
			if(en == 1) begin
				din[0]	<=	~key_1;
				din[1]	<=	din[0];
				if(din[0] == 1 && din[1] == 0) begin
					push	<=	1'b1;
				end
				else begin
					push	<=	1'b0;
				end
			end
			else begin
				din	<=	2'b0;
				push	<=	1'b0;
			end
		end
	end
	
	always @(posedge clk, negedge rstn) begin
		if(rstn == 0) begin
			rin	<=	2'd0;
			rpush	<=	1'b0;
		end
		else begin
			if(en == 1) begin
				rin[0]	<=	~iready;
				rin[1]	<=	rin[0];
				if(rin[0] == 1 && rin[1] == 0) begin
					rpush	<=	1'b1;
				end
				else begin
					rpush	<=	1'b0;
				end
			end
			else begin
				rin	<=	2'b0;
				rpush	<=	1'b0;
			end
		end
	end

	always @(posedge clk)
		if (rstn == 0)			cnt_en <= 0;
		else if (rpush)			cnt_en <= 1;
		else if (end_cnt_en)		cnt_en <= 0;

	always @(posedge clk)
		if (rstn == 0)	cnt <= 0;
		else if(cnt_en)	cnt <= cnt_max? 0: cnt + 1;

	always @(posedge clk)
		if (rstn == 0)	ready <= 0;
		else 		ready <= cnt_en;

	always @(posedge clk) begin
		if (cnt_en == 1'b0) begin
			dt	<=	1'b0;
		end
		else	begin
			case	(io)
				5'd2	:	begin
					case (cnt)
						10'd0	:	dt	<=	197	;
						10'd1	:	dt	<=	197	;
						10'd2	:	dt	<=	197	;
						10'd3	:	dt	<=	198	;
						10'd4	:	dt	<=	199	;
						10'd5	:	dt	<=	199	;
						10'd6	:	dt	<=	199	;
						10'd7	:	dt	<=	198	;
						10'd8	:	dt	<=	199	;
						10'd9	:	dt	<=	198	;
						10'd10	:	dt	<=	198	;
						10'd11	:	dt	<=	198	;
						10'd12	:	dt	<=	198	;
						10'd13	:	dt	<=	198	;
						10'd14	:	dt	<=	198	;
						10'd15	:	dt	<=	198	;
						10'd16	:	dt	<=	197	;
						10'd17	:	dt	<=	197	;
						10'd18	:	dt	<=	197	;
						10'd19	:	dt	<=	196	;
						10'd20	:	dt	<=	195	;
						10'd21	:	dt	<=	193	;
						10'd22	:	dt	<=	193	;
						10'd23	:	dt	<=	195	;
						10'd24	:	dt	<=	191	;
						10'd25	:	dt	<=	114	;
						10'd26	:	dt	<=	83	;
						10'd27	:	dt	<=	102	;
						10'd28	:	dt	<=	200	;
						10'd29	:	dt	<=	201	;
						10'd30	:	dt	<=	202	;
						10'd31	:	dt	<=	200	;
						10'd32	:	dt	<=	200	;
						10'd33	:	dt	<=	201	;
						10'd34	:	dt	<=	200	;
						10'd35	:	dt	<=	201	;
						10'd36	:	dt	<=	201	;
						10'd37	:	dt	<=	202	;
						10'd38	:	dt	<=	202	;
						10'd39	:	dt	<=	203	;
						10'd40	:	dt	<=	201	;
						10'd41	:	dt	<=	200	;
						10'd42	:	dt	<=	201	;
						10'd43	:	dt	<=	200	;
						10'd44	:	dt	<=	197	;
						10'd45	:	dt	<=	202	;
						10'd46	:	dt	<=	199	;
						10'd47	:	dt	<=	201	;
						10'd48	:	dt	<=	195	;
						10'd49	:	dt	<=	196	;
						10'd50	:	dt	<=	197	;
						10'd51	:	dt	<=	201	;
						10'd52	:	dt	<=	181	;
						10'd53	:	dt	<=	98	;
						10'd54	:	dt	<=	96	;
						10'd55	:	dt	<=	106	;
						10'd56	:	dt	<=	204	;
						10'd57	:	dt	<=	205	;
						10'd58	:	dt	<=	206	;
						10'd59	:	dt	<=	204	;
						10'd60	:	dt	<=	204	;
						10'd61	:	dt	<=	205	;
						10'd62	:	dt	<=	205	;
						10'd63	:	dt	<=	205	;
						10'd64	:	dt	<=	205	;
						10'd65	:	dt	<=	206	;
						10'd66	:	dt	<=	206	;
						10'd67	:	dt	<=	205	;
						10'd68	:	dt	<=	201	;
						10'd69	:	dt	<=	207	;
						10'd70	:	dt	<=	213	;
						10'd71	:	dt	<=	183	;
						10'd72	:	dt	<=	136	;
						10'd73	:	dt	<=	171	;
						10'd74	:	dt	<=	186	;
						10'd75	:	dt	<=	172	;
						10'd76	:	dt	<=	206	;
						10'd77	:	dt	<=	201	;
						10'd78	:	dt	<=	199	;
						10'd79	:	dt	<=	201	;
						10'd80	:	dt	<=	194	;
						10'd81	:	dt	<=	118	;
						10'd82	:	dt	<=	105	;
						10'd83	:	dt	<=	101	;
						10'd84	:	dt	<=	207	;
						10'd85	:	dt	<=	207	;
						10'd86	:	dt	<=	208	;
						10'd87	:	dt	<=	207	;
						10'd88	:	dt	<=	206	;
						10'd89	:	dt	<=	208	;
						10'd90	:	dt	<=	207	;
						10'd91	:	dt	<=	208	;
						10'd92	:	dt	<=	209	;
						10'd93	:	dt	<=	207	;
						10'd94	:	dt	<=	205	;
						10'd95	:	dt	<=	208	;
						10'd96	:	dt	<=	216	;
						10'd97	:	dt	<=	212	;
						10'd98	:	dt	<=	176	;
						10'd99	:	dt	<=	139	;
						10'd100	:	dt	<=	112	;
						10'd101	:	dt	<=	118	;
						10'd102	:	dt	<=	141	;
						10'd103	:	dt	<=	116	;
						10'd104	:	dt	<=	159	;
						10'd105	:	dt	<=	197	;
						10'd106	:	dt	<=	202	;
						10'd107	:	dt	<=	200	;
						10'd108	:	dt	<=	205	;
						10'd109	:	dt	<=	144	;
						10'd110	:	dt	<=	104	;
						10'd111	:	dt	<=	108	;
						10'd112	:	dt	<=	210	;
						10'd113	:	dt	<=	210	;
						10'd114	:	dt	<=	210	;
						10'd115	:	dt	<=	209	;
						10'd116	:	dt	<=	209	;
						10'd117	:	dt	<=	210	;
						10'd118	:	dt	<=	209	;
						10'd119	:	dt	<=	211	;
						10'd120	:	dt	<=	210	;
						10'd121	:	dt	<=	210	;
						10'd122	:	dt	<=	222	;
						10'd123	:	dt	<=	230	;
						10'd124	:	dt	<=	196	;
						10'd125	:	dt	<=	146	;
						10'd126	:	dt	<=	122	;
						10'd127	:	dt	<=	111	;
						10'd128	:	dt	<=	106	;
						10'd129	:	dt	<=	107	;
						10'd130	:	dt	<=	115	;
						10'd131	:	dt	<=	106	;
						10'd132	:	dt	<=	99	;
						10'd133	:	dt	<=	168	;
						10'd134	:	dt	<=	210	;
						10'd135	:	dt	<=	200	;
						10'd136	:	dt	<=	210	;
						10'd137	:	dt	<=	160	;
						10'd138	:	dt	<=	100	;
						10'd139	:	dt	<=	98	;
						10'd140	:	dt	<=	213	;
						10'd141	:	dt	<=	213	;
						10'd142	:	dt	<=	213	;
						10'd143	:	dt	<=	212	;
						10'd144	:	dt	<=	212	;
						10'd145	:	dt	<=	213	;
						10'd146	:	dt	<=	213	;
						10'd147	:	dt	<=	214	;
						10'd148	:	dt	<=	210	;
						10'd149	:	dt	<=	221	;
						10'd150	:	dt	<=	234	;
						10'd151	:	dt	<=	212	;
						10'd152	:	dt	<=	142	;
						10'd153	:	dt	<=	102	;
						10'd154	:	dt	<=	106	;
						10'd155	:	dt	<=	103	;
						10'd156	:	dt	<=	98	;
						10'd157	:	dt	<=	93	;
						10'd158	:	dt	<=	103	;
						10'd159	:	dt	<=	105	;
						10'd160	:	dt	<=	95	;
						10'd161	:	dt	<=	166	;
						10'd162	:	dt	<=	213	;
						10'd163	:	dt	<=	203	;
						10'd164	:	dt	<=	209	;
						10'd165	:	dt	<=	182	;
						10'd166	:	dt	<=	106	;
						10'd167	:	dt	<=	83	;
						10'd168	:	dt	<=	215	;
						10'd169	:	dt	<=	215	;
						10'd170	:	dt	<=	216	;
						10'd171	:	dt	<=	215	;
						10'd172	:	dt	<=	215	;
						10'd173	:	dt	<=	215	;
						10'd174	:	dt	<=	216	;
						10'd175	:	dt	<=	216	;
						10'd176	:	dt	<=	212	;
						10'd177	:	dt	<=	238	;
						10'd178	:	dt	<=	214	;
						10'd179	:	dt	<=	147	;
						10'd180	:	dt	<=	112	;
						10'd181	:	dt	<=	94	;
						10'd182	:	dt	<=	97	;
						10'd183	:	dt	<=	102	;
						10'd184	:	dt	<=	95	;
						10'd185	:	dt	<=	91	;
						10'd186	:	dt	<=	94	;
						10'd187	:	dt	<=	101	;
						10'd188	:	dt	<=	134	;
						10'd189	:	dt	<=	204	;
						10'd190	:	dt	<=	209	;
						10'd191	:	dt	<=	206	;
						10'd192	:	dt	<=	206	;
						10'd193	:	dt	<=	207	;
						10'd194	:	dt	<=	111	;
						10'd195	:	dt	<=	69	;
						10'd196	:	dt	<=	218	;
						10'd197	:	dt	<=	217	;
						10'd198	:	dt	<=	218	;
						10'd199	:	dt	<=	218	;
						10'd200	:	dt	<=	218	;
						10'd201	:	dt	<=	217	;
						10'd202	:	dt	<=	218	;
						10'd203	:	dt	<=	216	;
						10'd204	:	dt	<=	223	;
						10'd205	:	dt	<=	246	;
						10'd206	:	dt	<=	175	;
						10'd207	:	dt	<=	113	;
						10'd208	:	dt	<=	104	;
						10'd209	:	dt	<=	97	;
						10'd210	:	dt	<=	91	;
						10'd211	:	dt	<=	97	;
						10'd212	:	dt	<=	101	;
						10'd213	:	dt	<=	112	;
						10'd214	:	dt	<=	153	;
						10'd215	:	dt	<=	185	;
						10'd216	:	dt	<=	212	;
						10'd217	:	dt	<=	213	;
						10'd218	:	dt	<=	210	;
						10'd219	:	dt	<=	208	;
						10'd220	:	dt	<=	208	;
						10'd221	:	dt	<=	209	;
						10'd222	:	dt	<=	148	;
						10'd223	:	dt	<=	133	;
						10'd224	:	dt	<=	219	;
						10'd225	:	dt	<=	219	;
						10'd226	:	dt	<=	220	;
						10'd227	:	dt	<=	221	;
						10'd228	:	dt	<=	220	;
						10'd229	:	dt	<=	220	;
						10'd230	:	dt	<=	220	;
						10'd231	:	dt	<=	214	;
						10'd232	:	dt	<=	237	;
						10'd233	:	dt	<=	232	;
						10'd234	:	dt	<=	160	;
						10'd235	:	dt	<=	119	;
						10'd236	:	dt	<=	105	;
						10'd237	:	dt	<=	112	;
						10'd238	:	dt	<=	101	;
						10'd239	:	dt	<=	103	;
						10'd240	:	dt	<=	113	;
						10'd241	:	dt	<=	182	;
						10'd242	:	dt	<=	224	;
						10'd243	:	dt	<=	217	;
						10'd244	:	dt	<=	214	;
						10'd245	:	dt	<=	214	;
						10'd246	:	dt	<=	213	;
						10'd247	:	dt	<=	211	;
						10'd248	:	dt	<=	211	;
						10'd249	:	dt	<=	213	;
						10'd250	:	dt	<=	181	;
						10'd251	:	dt	<=	166	;
						10'd252	:	dt	<=	219	;
						10'd253	:	dt	<=	221	;
						10'd254	:	dt	<=	223	;
						10'd255	:	dt	<=	223	;
						10'd256	:	dt	<=	223	;
						10'd257	:	dt	<=	223	;
						10'd258	:	dt	<=	221	;
						10'd259	:	dt	<=	224	;
						10'd260	:	dt	<=	243	;
						10'd261	:	dt	<=	206	;
						10'd262	:	dt	<=	142	;
						10'd263	:	dt	<=	105	;
						10'd264	:	dt	<=	102	;
						10'd265	:	dt	<=	108	;
						10'd266	:	dt	<=	101	;
						10'd267	:	dt	<=	124	;
						10'd268	:	dt	<=	199	;
						10'd269	:	dt	<=	221	;
						10'd270	:	dt	<=	215	;
						10'd271	:	dt	<=	216	;
						10'd272	:	dt	<=	217	;
						10'd273	:	dt	<=	217	;
						10'd274	:	dt	<=	215	;
						10'd275	:	dt	<=	213	;
						10'd276	:	dt	<=	212	;
						10'd277	:	dt	<=	222	;
						10'd278	:	dt	<=	147	;
						10'd279	:	dt	<=	176	;
						10'd280	:	dt	<=	223	;
						10'd281	:	dt	<=	223	;
						10'd282	:	dt	<=	224	;
						10'd283	:	dt	<=	224	;
						10'd284	:	dt	<=	224	;
						10'd285	:	dt	<=	225	;
						10'd286	:	dt	<=	219	;
						10'd287	:	dt	<=	237	;
						10'd288	:	dt	<=	239	;
						10'd289	:	dt	<=	191	;
						10'd290	:	dt	<=	141	;
						10'd291	:	dt	<=	109	;
						10'd292	:	dt	<=	104	;
						10'd293	:	dt	<=	100	;
						10'd294	:	dt	<=	106	;
						10'd295	:	dt	<=	161	;
						10'd296	:	dt	<=	236	;
						10'd297	:	dt	<=	218	;
						10'd298	:	dt	<=	220	;
						10'd299	:	dt	<=	219	;
						10'd300	:	dt	<=	218	;
						10'd301	:	dt	<=	218	;
						10'd302	:	dt	<=	218	;
						10'd303	:	dt	<=	217	;
						10'd304	:	dt	<=	214	;
						10'd305	:	dt	<=	220	;
						10'd306	:	dt	<=	161	;
						10'd307	:	dt	<=	206	;
						10'd308	:	dt	<=	224	;
						10'd309	:	dt	<=	226	;
						10'd310	:	dt	<=	227	;
						10'd311	:	dt	<=	226	;
						10'd312	:	dt	<=	225	;
						10'd313	:	dt	<=	226	;
						10'd314	:	dt	<=	224	;
						10'd315	:	dt	<=	250	;
						10'd316	:	dt	<=	231	;
						10'd317	:	dt	<=	183	;
						10'd318	:	dt	<=	142	;
						10'd319	:	dt	<=	125	;
						10'd320	:	dt	<=	116	;
						10'd321	:	dt	<=	105	;
						10'd322	:	dt	<=	104	;
						10'd323	:	dt	<=	181	;
						10'd324	:	dt	<=	231	;
						10'd325	:	dt	<=	224	;
						10'd326	:	dt	<=	224	;
						10'd327	:	dt	<=	221	;
						10'd328	:	dt	<=	221	;
						10'd329	:	dt	<=	220	;
						10'd330	:	dt	<=	219	;
						10'd331	:	dt	<=	218	;
						10'd332	:	dt	<=	217	;
						10'd333	:	dt	<=	217	;
						10'd334	:	dt	<=	202	;
						10'd335	:	dt	<=	188	;
						10'd336	:	dt	<=	225	;
						10'd337	:	dt	<=	226	;
						10'd338	:	dt	<=	228	;
						10'd339	:	dt	<=	229	;
						10'd340	:	dt	<=	228	;
						10'd341	:	dt	<=	224	;
						10'd342	:	dt	<=	235	;
						10'd343	:	dt	<=	255	;
						10'd344	:	dt	<=	218	;
						10'd345	:	dt	<=	170	;
						10'd346	:	dt	<=	134	;
						10'd347	:	dt	<=	122	;
						10'd348	:	dt	<=	120	;
						10'd349	:	dt	<=	117	;
						10'd350	:	dt	<=	111	;
						10'd351	:	dt	<=	215	;
						10'd352	:	dt	<=	230	;
						10'd353	:	dt	<=	225	;
						10'd354	:	dt	<=	225	;
						10'd355	:	dt	<=	224	;
						10'd356	:	dt	<=	224	;
						10'd357	:	dt	<=	223	;
						10'd358	:	dt	<=	222	;
						10'd359	:	dt	<=	220	;
						10'd360	:	dt	<=	218	;
						10'd361	:	dt	<=	218	;
						10'd362	:	dt	<=	221	;
						10'd363	:	dt	<=	195	;
						10'd364	:	dt	<=	227	;
						10'd365	:	dt	<=	227	;
						10'd366	:	dt	<=	229	;
						10'd367	:	dt	<=	230	;
						10'd368	:	dt	<=	230	;
						10'd369	:	dt	<=	223	;
						10'd370	:	dt	<=	246	;
						10'd371	:	dt	<=	253	;
						10'd372	:	dt	<=	208	;
						10'd373	:	dt	<=	159	;
						10'd374	:	dt	<=	125	;
						10'd375	:	dt	<=	118	;
						10'd376	:	dt	<=	114	;
						10'd377	:	dt	<=	117	;
						10'd378	:	dt	<=	132	;
						10'd379	:	dt	<=	230	;
						10'd380	:	dt	<=	228	;
						10'd381	:	dt	<=	227	;
						10'd382	:	dt	<=	226	;
						10'd383	:	dt	<=	225	;
						10'd384	:	dt	<=	225	;
						10'd385	:	dt	<=	225	;
						10'd386	:	dt	<=	224	;
						10'd387	:	dt	<=	223	;
						10'd388	:	dt	<=	221	;
						10'd389	:	dt	<=	222	;
						10'd390	:	dt	<=	219	;
						10'd391	:	dt	<=	214	;
						10'd392	:	dt	<=	229	;
						10'd393	:	dt	<=	230	;
						10'd394	:	dt	<=	229	;
						10'd395	:	dt	<=	229	;
						10'd396	:	dt	<=	227	;
						10'd397	:	dt	<=	224	;
						10'd398	:	dt	<=	255	;
						10'd399	:	dt	<=	241	;
						10'd400	:	dt	<=	201	;
						10'd401	:	dt	<=	158	;
						10'd402	:	dt	<=	126	;
						10'd403	:	dt	<=	115	;
						10'd404	:	dt	<=	113	;
						10'd405	:	dt	<=	114	;
						10'd406	:	dt	<=	140	;
						10'd407	:	dt	<=	234	;
						10'd408	:	dt	<=	228	;
						10'd409	:	dt	<=	227	;
						10'd410	:	dt	<=	226	;
						10'd411	:	dt	<=	226	;
						10'd412	:	dt	<=	225	;
						10'd413	:	dt	<=	225	;
						10'd414	:	dt	<=	224	;
						10'd415	:	dt	<=	224	;
						10'd416	:	dt	<=	223	;
						10'd417	:	dt	<=	223	;
						10'd418	:	dt	<=	220	;
						10'd419	:	dt	<=	214	;
						10'd420	:	dt	<=	229	;
						10'd421	:	dt	<=	230	;
						10'd422	:	dt	<=	230	;
						10'd423	:	dt	<=	232	;
						10'd424	:	dt	<=	225	;
						10'd425	:	dt	<=	240	;
						10'd426	:	dt	<=	255	;
						10'd427	:	dt	<=	228	;
						10'd428	:	dt	<=	190	;
						10'd429	:	dt	<=	149	;
						10'd430	:	dt	<=	126	;
						10'd431	:	dt	<=	117	;
						10'd432	:	dt	<=	120	;
						10'd433	:	dt	<=	109	;
						10'd434	:	dt	<=	158	;
						10'd435	:	dt	<=	241	;
						10'd436	:	dt	<=	228	;
						10'd437	:	dt	<=	228	;
						10'd438	:	dt	<=	228	;
						10'd439	:	dt	<=	227	;
						10'd440	:	dt	<=	227	;
						10'd441	:	dt	<=	226	;
						10'd442	:	dt	<=	227	;
						10'd443	:	dt	<=	227	;
						10'd444	:	dt	<=	227	;
						10'd445	:	dt	<=	228	;
						10'd446	:	dt	<=	227	;
						10'd447	:	dt	<=	221	;
						10'd448	:	dt	<=	231	;
						10'd449	:	dt	<=	231	;
						10'd450	:	dt	<=	232	;
						10'd451	:	dt	<=	233	;
						10'd452	:	dt	<=	227	;
						10'd453	:	dt	<=	255	;
						10'd454	:	dt	<=	249	;
						10'd455	:	dt	<=	217	;
						10'd456	:	dt	<=	179	;
						10'd457	:	dt	<=	143	;
						10'd458	:	dt	<=	125	;
						10'd459	:	dt	<=	115	;
						10'd460	:	dt	<=	113	;
						10'd461	:	dt	<=	103	;
						10'd462	:	dt	<=	146	;
						10'd463	:	dt	<=	241	;
						10'd464	:	dt	<=	229	;
						10'd465	:	dt	<=	230	;
						10'd466	:	dt	<=	230	;
						10'd467	:	dt	<=	230	;
						10'd468	:	dt	<=	232	;
						10'd469	:	dt	<=	232	;
						10'd470	:	dt	<=	226	;
						10'd471	:	dt	<=	216	;
						10'd472	:	dt	<=	209	;
						10'd473	:	dt	<=	202	;
						10'd474	:	dt	<=	211	;
						10'd475	:	dt	<=	228	;
						10'd476	:	dt	<=	233	;
						10'd477	:	dt	<=	233	;
						10'd478	:	dt	<=	235	;
						10'd479	:	dt	<=	228	;
						10'd480	:	dt	<=	230	;
						10'd481	:	dt	<=	255	;
						10'd482	:	dt	<=	242	;
						10'd483	:	dt	<=	209	;
						10'd484	:	dt	<=	171	;
						10'd485	:	dt	<=	137	;
						10'd486	:	dt	<=	121	;
						10'd487	:	dt	<=	110	;
						10'd488	:	dt	<=	107	;
						10'd489	:	dt	<=	118	;
						10'd490	:	dt	<=	110	;
						10'd491	:	dt	<=	177	;
						10'd492	:	dt	<=	244	;
						10'd493	:	dt	<=	231	;
						10'd494	:	dt	<=	236	;
						10'd495	:	dt	<=	234	;
						10'd496	:	dt	<=	218	;
						10'd497	:	dt	<=	205	;
						10'd498	:	dt	<=	196	;
						10'd499	:	dt	<=	193	;
						10'd500	:	dt	<=	189	;
						10'd501	:	dt	<=	178	;
						10'd502	:	dt	<=	151	;
						10'd503	:	dt	<=	181	;
						10'd504	:	dt	<=	233	;
						10'd505	:	dt	<=	234	;
						10'd506	:	dt	<=	238	;
						10'd507	:	dt	<=	224	;
						10'd508	:	dt	<=	243	;
						10'd509	:	dt	<=	255	;
						10'd510	:	dt	<=	235	;
						10'd511	:	dt	<=	199	;
						10'd512	:	dt	<=	162	;
						10'd513	:	dt	<=	136	;
						10'd514	:	dt	<=	118	;
						10'd515	:	dt	<=	100	;
						10'd516	:	dt	<=	110	;
						10'd517	:	dt	<=	121	;
						10'd518	:	dt	<=	123	;
						10'd519	:	dt	<=	117	;
						10'd520	:	dt	<=	207	;
						10'd521	:	dt	<=	233	;
						10'd522	:	dt	<=	218	;
						10'd523	:	dt	<=	198	;
						10'd524	:	dt	<=	191	;
						10'd525	:	dt	<=	192	;
						10'd526	:	dt	<=	202	;
						10'd527	:	dt	<=	196	;
						10'd528	:	dt	<=	175	;
						10'd529	:	dt	<=	158	;
						10'd530	:	dt	<=	146	;
						10'd531	:	dt	<=	166	;
						10'd532	:	dt	<=	235	;
						10'd533	:	dt	<=	237	;
						10'd534	:	dt	<=	233	;
						10'd535	:	dt	<=	229	;
						10'd536	:	dt	<=	255	;
						10'd537	:	dt	<=	251	;
						10'd538	:	dt	<=	225	;
						10'd539	:	dt	<=	185	;
						10'd540	:	dt	<=	152	;
						10'd541	:	dt	<=	134	;
						10'd542	:	dt	<=	111	;
						10'd543	:	dt	<=	96	;
						10'd544	:	dt	<=	118	;
						10'd545	:	dt	<=	122	;
						10'd546	:	dt	<=	128	;
						10'd547	:	dt	<=	135	;
						10'd548	:	dt	<=	136	;
						10'd549	:	dt	<=	159	;
						10'd550	:	dt	<=	172	;
						10'd551	:	dt	<=	190	;
						10'd552	:	dt	<=	205	;
						10'd553	:	dt	<=	197	;
						10'd554	:	dt	<=	177	;
						10'd555	:	dt	<=	146	;
						10'd556	:	dt	<=	154	;
						10'd557	:	dt	<=	200	;
						10'd558	:	dt	<=	222	;
						10'd559	:	dt	<=	228	;
						10'd560	:	dt	<=	237	;
						10'd561	:	dt	<=	240	;
						10'd562	:	dt	<=	227	;
						10'd563	:	dt	<=	244	;
						10'd564	:	dt	<=	255	;
						10'd565	:	dt	<=	243	;
						10'd566	:	dt	<=	216	;
						10'd567	:	dt	<=	178	;
						10'd568	:	dt	<=	149	;
						10'd569	:	dt	<=	131	;
						10'd570	:	dt	<=	104	;
						10'd571	:	dt	<=	106	;
						10'd572	:	dt	<=	132	;
						10'd573	:	dt	<=	136	;
						10'd574	:	dt	<=	147	;
						10'd575	:	dt	<=	149	;
						10'd576	:	dt	<=	147	;
						10'd577	:	dt	<=	154	;
						10'd578	:	dt	<=	178	;
						10'd579	:	dt	<=	196	;
						10'd580	:	dt	<=	185	;
						10'd581	:	dt	<=	155	;
						10'd582	:	dt	<=	129	;
						10'd583	:	dt	<=	160	;
						10'd584	:	dt	<=	229	;
						10'd585	:	dt	<=	234	;
						10'd586	:	dt	<=	232	;
						10'd587	:	dt	<=	231	;
						10'd588	:	dt	<=	240	;
						10'd589	:	dt	<=	234	;
						10'd590	:	dt	<=	231	;
						10'd591	:	dt	<=	255	;
						10'd592	:	dt	<=	253	;
						10'd593	:	dt	<=	237	;
						10'd594	:	dt	<=	204	;
						10'd595	:	dt	<=	172	;
						10'd596	:	dt	<=	146	;
						10'd597	:	dt	<=	130	;
						10'd598	:	dt	<=	105	;
						10'd599	:	dt	<=	118	;
						10'd600	:	dt	<=	142	;
						10'd601	:	dt	<=	149	;
						10'd602	:	dt	<=	154	;
						10'd603	:	dt	<=	151	;
						10'd604	:	dt	<=	152	;
						10'd605	:	dt	<=	157	;
						10'd606	:	dt	<=	168	;
						10'd607	:	dt	<=	152	;
						10'd608	:	dt	<=	144	;
						10'd609	:	dt	<=	166	;
						10'd610	:	dt	<=	199	;
						10'd611	:	dt	<=	234	;
						10'd612	:	dt	<=	234	;
						10'd613	:	dt	<=	230	;
						10'd614	:	dt	<=	230	;
						10'd615	:	dt	<=	229	;
						10'd616	:	dt	<=	237	;
						10'd617	:	dt	<=	230	;
						10'd618	:	dt	<=	253	;
						10'd619	:	dt	<=	255	;
						10'd620	:	dt	<=	246	;
						10'd621	:	dt	<=	228	;
						10'd622	:	dt	<=	198	;
						10'd623	:	dt	<=	165	;
						10'd624	:	dt	<=	136	;
						10'd625	:	dt	<=	127	;
						10'd626	:	dt	<=	112	;
						10'd627	:	dt	<=	129	;
						10'd628	:	dt	<=	147	;
						10'd629	:	dt	<=	156	;
						10'd630	:	dt	<=	157	;
						10'd631	:	dt	<=	152	;
						10'd632	:	dt	<=	144	;
						10'd633	:	dt	<=	136	;
						10'd634	:	dt	<=	130	;
						10'd635	:	dt	<=	160	;
						10'd636	:	dt	<=	213	;
						10'd637	:	dt	<=	239	;
						10'd638	:	dt	<=	240	;
						10'd639	:	dt	<=	235	;
						10'd640	:	dt	<=	234	;
						10'd641	:	dt	<=	233	;
						10'd642	:	dt	<=	232	;
						10'd643	:	dt	<=	231	;
						10'd644	:	dt	<=	225	;
						10'd645	:	dt	<=	242	;
						10'd646	:	dt	<=	255	;
						10'd647	:	dt	<=	249	;
						10'd648	:	dt	<=	241	;
						10'd649	:	dt	<=	225	;
						10'd650	:	dt	<=	191	;
						10'd651	:	dt	<=	156	;
						10'd652	:	dt	<=	131	;
						10'd653	:	dt	<=	127	;
						10'd654	:	dt	<=	119	;
						10'd655	:	dt	<=	142	;
						10'd656	:	dt	<=	153	;
						10'd657	:	dt	<=	155	;
						10'd658	:	dt	<=	150	;
						10'd659	:	dt	<=	139	;
						10'd660	:	dt	<=	125	;
						10'd661	:	dt	<=	131	;
						10'd662	:	dt	<=	189	;
						10'd663	:	dt	<=	241	;
						10'd664	:	dt	<=	241	;
						10'd665	:	dt	<=	237	;
						10'd666	:	dt	<=	236	;
						10'd667	:	dt	<=	236	;
						10'd668	:	dt	<=	236	;
						10'd669	:	dt	<=	235	;
						10'd670	:	dt	<=	235	;
						10'd671	:	dt	<=	234	;
						10'd672	:	dt	<=	236	;
						10'd673	:	dt	<=	247	;
						10'd674	:	dt	<=	248	;
						10'd675	:	dt	<=	241	;
						10'd676	:	dt	<=	229	;
						10'd677	:	dt	<=	203	;
						10'd678	:	dt	<=	169	;
						10'd679	:	dt	<=	142	;
						10'd680	:	dt	<=	131	;
						10'd681	:	dt	<=	123	;
						10'd682	:	dt	<=	126	;
						10'd683	:	dt	<=	145	;
						10'd684	:	dt	<=	148	;
						10'd685	:	dt	<=	150	;
						10'd686	:	dt	<=	135	;
						10'd687	:	dt	<=	122	;
						10'd688	:	dt	<=	172	;
						10'd689	:	dt	<=	224	;
						10'd690	:	dt	<=	245	;
						10'd691	:	dt	<=	239	;
						10'd692	:	dt	<=	238	;
						10'd693	:	dt	<=	240	;
						10'd694	:	dt	<=	239	;
						10'd695	:	dt	<=	238	;
						10'd696	:	dt	<=	237	;
						10'd697	:	dt	<=	236	;
						10'd698	:	dt	<=	236	;
						10'd699	:	dt	<=	236	;
						10'd700	:	dt	<=	243	;
						10'd701	:	dt	<=	245	;
						10'd702	:	dt	<=	240	;
						10'd703	:	dt	<=	222	;
						10'd704	:	dt	<=	202	;
						10'd705	:	dt	<=	177	;
						10'd706	:	dt	<=	153	;
						10'd707	:	dt	<=	135	;
						10'd708	:	dt	<=	130	;
						10'd709	:	dt	<=	124	;
						10'd710	:	dt	<=	132	;
						10'd711	:	dt	<=	138	;
						10'd712	:	dt	<=	143	;
						10'd713	:	dt	<=	136	;
						10'd714	:	dt	<=	120	;
						10'd715	:	dt	<=	187	;
						10'd716	:	dt	<=	249	;
						10'd717	:	dt	<=	245	;
						10'd718	:	dt	<=	239	;
						10'd719	:	dt	<=	240	;
						10'd720	:	dt	<=	240	;
						10'd721	:	dt	<=	241	;
						10'd722	:	dt	<=	241	;
						10'd723	:	dt	<=	241	;
						10'd724	:	dt	<=	239	;
						10'd725	:	dt	<=	238	;
						10'd726	:	dt	<=	238	;
						10'd727	:	dt	<=	237	;
						10'd728	:	dt	<=	240	;
						10'd729	:	dt	<=	239	;
						10'd730	:	dt	<=	224	;
						10'd731	:	dt	<=	202	;
						10'd732	:	dt	<=	184	;
						10'd733	:	dt	<=	168	;
						10'd734	:	dt	<=	146	;
						10'd735	:	dt	<=	132	;
						10'd736	:	dt	<=	128	;
						10'd737	:	dt	<=	131	;
						10'd738	:	dt	<=	131	;
						10'd739	:	dt	<=	130	;
						10'd740	:	dt	<=	128	;
						10'd741	:	dt	<=	138	;
						10'd742	:	dt	<=	203	;
						10'd743	:	dt	<=	249	;
						10'd744	:	dt	<=	241	;
						10'd745	:	dt	<=	242	;
						10'd746	:	dt	<=	243	;
						10'd747	:	dt	<=	242	;
						10'd748	:	dt	<=	242	;
						10'd749	:	dt	<=	242	;
						10'd750	:	dt	<=	242	;
						10'd751	:	dt	<=	242	;
						10'd752	:	dt	<=	240	;
						10'd753	:	dt	<=	239	;
						10'd754	:	dt	<=	237	;
						10'd755	:	dt	<=	236	;
						10'd756	:	dt	<=	238	;
						10'd757	:	dt	<=	230	;
						10'd758	:	dt	<=	211	;
						10'd759	:	dt	<=	180	;
						10'd760	:	dt	<=	170	;
						10'd761	:	dt	<=	149	;
						10'd762	:	dt	<=	130	;
						10'd763	:	dt	<=	132	;
						10'd764	:	dt	<=	133	;
						10'd765	:	dt	<=	132	;
						10'd766	:	dt	<=	130	;
						10'd767	:	dt	<=	124	;
						10'd768	:	dt	<=	172	;
						10'd769	:	dt	<=	236	;
						10'd770	:	dt	<=	250	;
						10'd771	:	dt	<=	243	;
						10'd772	:	dt	<=	245	;
						10'd773	:	dt	<=	245	;
						10'd774	:	dt	<=	244	;
						10'd775	:	dt	<=	245	;
						10'd776	:	dt	<=	244	;
						10'd777	:	dt	<=	243	;
						10'd778	:	dt	<=	243	;
						10'd779	:	dt	<=	242	;
						10'd780	:	dt	<=	241	;
						10'd781	:	dt	<=	240	;
						10'd782	:	dt	<=	239	;
						10'd783	:	dt	<=	238	;
					endcase
				end
				5'd4	:	begin
					case (cnt)
						10'd0	:	dt	<=	191	;
						10'd1	:	dt	<=	192	;
						10'd2	:	dt	<=	192	;
						10'd3	:	dt	<=	192	;
						10'd4	:	dt	<=	192	;
						10'd5	:	dt	<=	193	;
						10'd6	:	dt	<=	193	;
						10'd7	:	dt	<=	193	;
						10'd8	:	dt	<=	193	;
						10'd9	:	dt	<=	192	;
						10'd10	:	dt	<=	193	;
						10'd11	:	dt	<=	193	;
						10'd12	:	dt	<=	192	;
						10'd13	:	dt	<=	192	;
						10'd14	:	dt	<=	192	;
						10'd15	:	dt	<=	191	;
						10'd16	:	dt	<=	190	;
						10'd17	:	dt	<=	187	;
						10'd18	:	dt	<=	188	;
						10'd19	:	dt	<=	188	;
						10'd20	:	dt	<=	187	;
						10'd21	:	dt	<=	186	;
						10'd22	:	dt	<=	184	;
						10'd23	:	dt	<=	184	;
						10'd24	:	dt	<=	182	;
						10'd25	:	dt	<=	182	;
						10'd26	:	dt	<=	181	;
						10'd27	:	dt	<=	180	;
						10'd28	:	dt	<=	193	;
						10'd29	:	dt	<=	194	;
						10'd30	:	dt	<=	195	;
						10'd31	:	dt	<=	195	;
						10'd32	:	dt	<=	195	;
						10'd33	:	dt	<=	195	;
						10'd34	:	dt	<=	195	;
						10'd35	:	dt	<=	195	;
						10'd36	:	dt	<=	195	;
						10'd37	:	dt	<=	194	;
						10'd38	:	dt	<=	194	;
						10'd39	:	dt	<=	195	;
						10'd40	:	dt	<=	196	;
						10'd41	:	dt	<=	194	;
						10'd42	:	dt	<=	193	;
						10'd43	:	dt	<=	193	;
						10'd44	:	dt	<=	193	;
						10'd45	:	dt	<=	195	;
						10'd46	:	dt	<=	192	;
						10'd47	:	dt	<=	189	;
						10'd48	:	dt	<=	188	;
						10'd49	:	dt	<=	187	;
						10'd50	:	dt	<=	187	;
						10'd51	:	dt	<=	186	;
						10'd52	:	dt	<=	185	;
						10'd53	:	dt	<=	184	;
						10'd54	:	dt	<=	183	;
						10'd55	:	dt	<=	181	;
						10'd56	:	dt	<=	198	;
						10'd57	:	dt	<=	197	;
						10'd58	:	dt	<=	198	;
						10'd59	:	dt	<=	197	;
						10'd60	:	dt	<=	197	;
						10'd61	:	dt	<=	198	;
						10'd62	:	dt	<=	197	;
						10'd63	:	dt	<=	197	;
						10'd64	:	dt	<=	197	;
						10'd65	:	dt	<=	198	;
						10'd66	:	dt	<=	197	;
						10'd67	:	dt	<=	195	;
						10'd68	:	dt	<=	193	;
						10'd69	:	dt	<=	199	;
						10'd70	:	dt	<=	198	;
						10'd71	:	dt	<=	189	;
						10'd72	:	dt	<=	164	;
						10'd73	:	dt	<=	155	;
						10'd74	:	dt	<=	190	;
						10'd75	:	dt	<=	195	;
						10'd76	:	dt	<=	194	;
						10'd77	:	dt	<=	193	;
						10'd78	:	dt	<=	188	;
						10'd79	:	dt	<=	188	;
						10'd80	:	dt	<=	188	;
						10'd81	:	dt	<=	187	;
						10'd82	:	dt	<=	186	;
						10'd83	:	dt	<=	185	;
						10'd84	:	dt	<=	200	;
						10'd85	:	dt	<=	199	;
						10'd86	:	dt	<=	199	;
						10'd87	:	dt	<=	200	;
						10'd88	:	dt	<=	199	;
						10'd89	:	dt	<=	199	;
						10'd90	:	dt	<=	199	;
						10'd91	:	dt	<=	199	;
						10'd92	:	dt	<=	199	;
						10'd93	:	dt	<=	198	;
						10'd94	:	dt	<=	197	;
						10'd95	:	dt	<=	183	;
						10'd96	:	dt	<=	159	;
						10'd97	:	dt	<=	161	;
						10'd98	:	dt	<=	197	;
						10'd99	:	dt	<=	192	;
						10'd100	:	dt	<=	163	;
						10'd101	:	dt	<=	122	;
						10'd102	:	dt	<=	145	;
						10'd103	:	dt	<=	193	;
						10'd104	:	dt	<=	159	;
						10'd105	:	dt	<=	168	;
						10'd106	:	dt	<=	193	;
						10'd107	:	dt	<=	190	;
						10'd108	:	dt	<=	189	;
						10'd109	:	dt	<=	189	;
						10'd110	:	dt	<=	187	;
						10'd111	:	dt	<=	186	;
						10'd112	:	dt	<=	202	;
						10'd113	:	dt	<=	201	;
						10'd114	:	dt	<=	201	;
						10'd115	:	dt	<=	202	;
						10'd116	:	dt	<=	202	;
						10'd117	:	dt	<=	201	;
						10'd118	:	dt	<=	201	;
						10'd119	:	dt	<=	201	;
						10'd120	:	dt	<=	201	;
						10'd121	:	dt	<=	200	;
						10'd122	:	dt	<=	204	;
						10'd123	:	dt	<=	207	;
						10'd124	:	dt	<=	182	;
						10'd125	:	dt	<=	152	;
						10'd126	:	dt	<=	141	;
						10'd127	:	dt	<=	187	;
						10'd128	:	dt	<=	181	;
						10'd129	:	dt	<=	145	;
						10'd130	:	dt	<=	108	;
						10'd131	:	dt	<=	159	;
						10'd132	:	dt	<=	152	;
						10'd133	:	dt	<=	111	;
						10'd134	:	dt	<=	157	;
						10'd135	:	dt	<=	200	;
						10'd136	:	dt	<=	189	;
						10'd137	:	dt	<=	191	;
						10'd138	:	dt	<=	189	;
						10'd139	:	dt	<=	188	;
						10'd140	:	dt	<=	202	;
						10'd141	:	dt	<=	202	;
						10'd142	:	dt	<=	203	;
						10'd143	:	dt	<=	204	;
						10'd144	:	dt	<=	204	;
						10'd145	:	dt	<=	203	;
						10'd146	:	dt	<=	203	;
						10'd147	:	dt	<=	204	;
						10'd148	:	dt	<=	202	;
						10'd149	:	dt	<=	196	;
						10'd150	:	dt	<=	193	;
						10'd151	:	dt	<=	196	;
						10'd152	:	dt	<=	203	;
						10'd153	:	dt	<=	181	;
						10'd154	:	dt	<=	136	;
						10'd155	:	dt	<=	136	;
						10'd156	:	dt	<=	186	;
						10'd157	:	dt	<=	163	;
						10'd158	:	dt	<=	110	;
						10'd159	:	dt	<=	136	;
						10'd160	:	dt	<=	162	;
						10'd161	:	dt	<=	116	;
						10'd162	:	dt	<=	107	;
						10'd163	:	dt	<=	198	;
						10'd164	:	dt	<=	192	;
						10'd165	:	dt	<=	193	;
						10'd166	:	dt	<=	191	;
						10'd167	:	dt	<=	190	;
						10'd168	:	dt	<=	205	;
						10'd169	:	dt	<=	204	;
						10'd170	:	dt	<=	204	;
						10'd171	:	dt	<=	205	;
						10'd172	:	dt	<=	205	;
						10'd173	:	dt	<=	206	;
						10'd174	:	dt	<=	205	;
						10'd175	:	dt	<=	207	;
						10'd176	:	dt	<=	198	;
						10'd177	:	dt	<=	187	;
						10'd178	:	dt	<=	185	;
						10'd179	:	dt	<=	143	;
						10'd180	:	dt	<=	163	;
						10'd181	:	dt	<=	180	;
						10'd182	:	dt	<=	123	;
						10'd183	:	dt	<=	105	;
						10'd184	:	dt	<=	183	;
						10'd185	:	dt	<=	162	;
						10'd186	:	dt	<=	110	;
						10'd187	:	dt	<=	117	;
						10'd188	:	dt	<=	164	;
						10'd189	:	dt	<=	131	;
						10'd190	:	dt	<=	95	;
						10'd191	:	dt	<=	193	;
						10'd192	:	dt	<=	195	;
						10'd193	:	dt	<=	193	;
						10'd194	:	dt	<=	192	;
						10'd195	:	dt	<=	191	;
						10'd196	:	dt	<=	206	;
						10'd197	:	dt	<=	206	;
						10'd198	:	dt	<=	207	;
						10'd199	:	dt	<=	207	;
						10'd200	:	dt	<=	207	;
						10'd201	:	dt	<=	206	;
						10'd202	:	dt	<=	207	;
						10'd203	:	dt	<=	206	;
						10'd204	:	dt	<=	201	;
						10'd205	:	dt	<=	198	;
						10'd206	:	dt	<=	189	;
						10'd207	:	dt	<=	142	;
						10'd208	:	dt	<=	120	;
						10'd209	:	dt	<=	161	;
						10'd210	:	dt	<=	115	;
						10'd211	:	dt	<=	99	;
						10'd212	:	dt	<=	164	;
						10'd213	:	dt	<=	133	;
						10'd214	:	dt	<=	90	;
						10'd215	:	dt	<=	137	;
						10'd216	:	dt	<=	169	;
						10'd217	:	dt	<=	137	;
						10'd218	:	dt	<=	107	;
						10'd219	:	dt	<=	200	;
						10'd220	:	dt	<=	197	;
						10'd221	:	dt	<=	196	;
						10'd222	:	dt	<=	195	;
						10'd223	:	dt	<=	195	;
						10'd224	:	dt	<=	207	;
						10'd225	:	dt	<=	207	;
						10'd226	:	dt	<=	208	;
						10'd227	:	dt	<=	207	;
						10'd228	:	dt	<=	208	;
						10'd229	:	dt	<=	208	;
						10'd230	:	dt	<=	208	;
						10'd231	:	dt	<=	209	;
						10'd232	:	dt	<=	194	;
						10'd233	:	dt	<=	154	;
						10'd234	:	dt	<=	181	;
						10'd235	:	dt	<=	158	;
						10'd236	:	dt	<=	114	;
						10'd237	:	dt	<=	141	;
						10'd238	:	dt	<=	146	;
						10'd239	:	dt	<=	97	;
						10'd240	:	dt	<=	133	;
						10'd241	:	dt	<=	120	;
						10'd242	:	dt	<=	78	;
						10'd243	:	dt	<=	144	;
						10'd244	:	dt	<=	143	;
						10'd245	:	dt	<=	102	;
						10'd246	:	dt	<=	123	;
						10'd247	:	dt	<=	209	;
						10'd248	:	dt	<=	197	;
						10'd249	:	dt	<=	198	;
						10'd250	:	dt	<=	198	;
						10'd251	:	dt	<=	196	;
						10'd252	:	dt	<=	209	;
						10'd253	:	dt	<=	208	;
						10'd254	:	dt	<=	209	;
						10'd255	:	dt	<=	209	;
						10'd256	:	dt	<=	209	;
						10'd257	:	dt	<=	209	;
						10'd258	:	dt	<=	209	;
						10'd259	:	dt	<=	208	;
						10'd260	:	dt	<=	207	;
						10'd261	:	dt	<=	154	;
						10'd262	:	dt	<=	140	;
						10'd263	:	dt	<=	182	;
						10'd264	:	dt	<=	144	;
						10'd265	:	dt	<=	124	;
						10'd266	:	dt	<=	172	;
						10'd267	:	dt	<=	105	;
						10'd268	:	dt	<=	112	;
						10'd269	:	dt	<=	137	;
						10'd270	:	dt	<=	133	;
						10'd271	:	dt	<=	138	;
						10'd272	:	dt	<=	105	;
						10'd273	:	dt	<=	68	;
						10'd274	:	dt	<=	145	;
						10'd275	:	dt	<=	212	;
						10'd276	:	dt	<=	199	;
						10'd277	:	dt	<=	200	;
						10'd278	:	dt	<=	199	;
						10'd279	:	dt	<=	198	;
						10'd280	:	dt	<=	210	;
						10'd281	:	dt	<=	210	;
						10'd282	:	dt	<=	209	;
						10'd283	:	dt	<=	210	;
						10'd284	:	dt	<=	211	;
						10'd285	:	dt	<=	209	;
						10'd286	:	dt	<=	208	;
						10'd287	:	dt	<=	211	;
						10'd288	:	dt	<=	196	;
						10'd289	:	dt	<=	138	;
						10'd290	:	dt	<=	113	;
						10'd291	:	dt	<=	172	;
						10'd292	:	dt	<=	148	;
						10'd293	:	dt	<=	164	;
						10'd294	:	dt	<=	171	;
						10'd295	:	dt	<=	151	;
						10'd296	:	dt	<=	154	;
						10'd297	:	dt	<=	153	;
						10'd298	:	dt	<=	179	;
						10'd299	:	dt	<=	150	;
						10'd300	:	dt	<=	94	;
						10'd301	:	dt	<=	72	;
						10'd302	:	dt	<=	182	;
						10'd303	:	dt	<=	207	;
						10'd304	:	dt	<=	201	;
						10'd305	:	dt	<=	202	;
						10'd306	:	dt	<=	200	;
						10'd307	:	dt	<=	199	;
						10'd308	:	dt	<=	210	;
						10'd309	:	dt	<=	210	;
						10'd310	:	dt	<=	211	;
						10'd311	:	dt	<=	211	;
						10'd312	:	dt	<=	210	;
						10'd313	:	dt	<=	210	;
						10'd314	:	dt	<=	210	;
						10'd315	:	dt	<=	212	;
						10'd316	:	dt	<=	196	;
						10'd317	:	dt	<=	171	;
						10'd318	:	dt	<=	168	;
						10'd319	:	dt	<=	140	;
						10'd320	:	dt	<=	94	;
						10'd321	:	dt	<=	181	;
						10'd322	:	dt	<=	171	;
						10'd323	:	dt	<=	160	;
						10'd324	:	dt	<=	169	;
						10'd325	:	dt	<=	157	;
						10'd326	:	dt	<=	167	;
						10'd327	:	dt	<=	141	;
						10'd328	:	dt	<=	102	;
						10'd329	:	dt	<=	95	;
						10'd330	:	dt	<=	206	;
						10'd331	:	dt	<=	204	;
						10'd332	:	dt	<=	203	;
						10'd333	:	dt	<=	203	;
						10'd334	:	dt	<=	202	;
						10'd335	:	dt	<=	200	;
						10'd336	:	dt	<=	211	;
						10'd337	:	dt	<=	211	;
						10'd338	:	dt	<=	211	;
						10'd339	:	dt	<=	211	;
						10'd340	:	dt	<=	212	;
						10'd341	:	dt	<=	212	;
						10'd342	:	dt	<=	211	;
						10'd343	:	dt	<=	211	;
						10'd344	:	dt	<=	207	;
						10'd345	:	dt	<=	193	;
						10'd346	:	dt	<=	156	;
						10'd347	:	dt	<=	120	;
						10'd348	:	dt	<=	88	;
						10'd349	:	dt	<=	117	;
						10'd350	:	dt	<=	148	;
						10'd351	:	dt	<=	137	;
						10'd352	:	dt	<=	140	;
						10'd353	:	dt	<=	137	;
						10'd354	:	dt	<=	131	;
						10'd355	:	dt	<=	130	;
						10'd356	:	dt	<=	120	;
						10'd357	:	dt	<=	93	;
						10'd358	:	dt	<=	179	;
						10'd359	:	dt	<=	213	;
						10'd360	:	dt	<=	204	;
						10'd361	:	dt	<=	204	;
						10'd362	:	dt	<=	203	;
						10'd363	:	dt	<=	201	;
						10'd364	:	dt	<=	212	;
						10'd365	:	dt	<=	212	;
						10'd366	:	dt	<=	212	;
						10'd367	:	dt	<=	212	;
						10'd368	:	dt	<=	213	;
						10'd369	:	dt	<=	212	;
						10'd370	:	dt	<=	211	;
						10'd371	:	dt	<=	210	;
						10'd372	:	dt	<=	208	;
						10'd373	:	dt	<=	181	;
						10'd374	:	dt	<=	142	;
						10'd375	:	dt	<=	109	;
						10'd376	:	dt	<=	99	;
						10'd377	:	dt	<=	97	;
						10'd378	:	dt	<=	115	;
						10'd379	:	dt	<=	125	;
						10'd380	:	dt	<=	125	;
						10'd381	:	dt	<=	120	;
						10'd382	:	dt	<=	112	;
						10'd383	:	dt	<=	141	;
						10'd384	:	dt	<=	135	;
						10'd385	:	dt	<=	108	;
						10'd386	:	dt	<=	110	;
						10'd387	:	dt	<=	211	;
						10'd388	:	dt	<=	206	;
						10'd389	:	dt	<=	205	;
						10'd390	:	dt	<=	205	;
						10'd391	:	dt	<=	204	;
						10'd392	:	dt	<=	213	;
						10'd393	:	dt	<=	213	;
						10'd394	:	dt	<=	213	;
						10'd395	:	dt	<=	213	;
						10'd396	:	dt	<=	213	;
						10'd397	:	dt	<=	214	;
						10'd398	:	dt	<=	212	;
						10'd399	:	dt	<=	210	;
						10'd400	:	dt	<=	200	;
						10'd401	:	dt	<=	164	;
						10'd402	:	dt	<=	130	;
						10'd403	:	dt	<=	106	;
						10'd404	:	dt	<=	103	;
						10'd405	:	dt	<=	122	;
						10'd406	:	dt	<=	127	;
						10'd407	:	dt	<=	155	;
						10'd408	:	dt	<=	164	;
						10'd409	:	dt	<=	159	;
						10'd410	:	dt	<=	141	;
						10'd411	:	dt	<=	148	;
						10'd412	:	dt	<=	149	;
						10'd413	:	dt	<=	140	;
						10'd414	:	dt	<=	92	;
						10'd415	:	dt	<=	160	;
						10'd416	:	dt	<=	217	;
						10'd417	:	dt	<=	203	;
						10'd418	:	dt	<=	205	;
						10'd419	:	dt	<=	204	;
						10'd420	:	dt	<=	214	;
						10'd421	:	dt	<=	215	;
						10'd422	:	dt	<=	215	;
						10'd423	:	dt	<=	215	;
						10'd424	:	dt	<=	215	;
						10'd425	:	dt	<=	215	;
						10'd426	:	dt	<=	213	;
						10'd427	:	dt	<=	207	;
						10'd428	:	dt	<=	201	;
						10'd429	:	dt	<=	175	;
						10'd430	:	dt	<=	143	;
						10'd431	:	dt	<=	113	;
						10'd432	:	dt	<=	115	;
						10'd433	:	dt	<=	122	;
						10'd434	:	dt	<=	146	;
						10'd435	:	dt	<=	183	;
						10'd436	:	dt	<=	183	;
						10'd437	:	dt	<=	197	;
						10'd438	:	dt	<=	184	;
						10'd439	:	dt	<=	159	;
						10'd440	:	dt	<=	186	;
						10'd441	:	dt	<=	161	;
						10'd442	:	dt	<=	109	;
						10'd443	:	dt	<=	106	;
						10'd444	:	dt	<=	214	;
						10'd445	:	dt	<=	206	;
						10'd446	:	dt	<=	206	;
						10'd447	:	dt	<=	205	;
						10'd448	:	dt	<=	216	;
						10'd449	:	dt	<=	216	;
						10'd450	:	dt	<=	215	;
						10'd451	:	dt	<=	216	;
						10'd452	:	dt	<=	216	;
						10'd453	:	dt	<=	216	;
						10'd454	:	dt	<=	215	;
						10'd455	:	dt	<=	205	;
						10'd456	:	dt	<=	202	;
						10'd457	:	dt	<=	178	;
						10'd458	:	dt	<=	144	;
						10'd459	:	dt	<=	111	;
						10'd460	:	dt	<=	111	;
						10'd461	:	dt	<=	131	;
						10'd462	:	dt	<=	164	;
						10'd463	:	dt	<=	193	;
						10'd464	:	dt	<=	194	;
						10'd465	:	dt	<=	205	;
						10'd466	:	dt	<=	209	;
						10'd467	:	dt	<=	191	;
						10'd468	:	dt	<=	175	;
						10'd469	:	dt	<=	160	;
						10'd470	:	dt	<=	106	;
						10'd471	:	dt	<=	101	;
						10'd472	:	dt	<=	213	;
						10'd473	:	dt	<=	208	;
						10'd474	:	dt	<=	207	;
						10'd475	:	dt	<=	206	;
						10'd476	:	dt	<=	216	;
						10'd477	:	dt	<=	217	;
						10'd478	:	dt	<=	216	;
						10'd479	:	dt	<=	216	;
						10'd480	:	dt	<=	216	;
						10'd481	:	dt	<=	217	;
						10'd482	:	dt	<=	216	;
						10'd483	:	dt	<=	199	;
						10'd484	:	dt	<=	200	;
						10'd485	:	dt	<=	188	;
						10'd486	:	dt	<=	152	;
						10'd487	:	dt	<=	119	;
						10'd488	:	dt	<=	117	;
						10'd489	:	dt	<=	133	;
						10'd490	:	dt	<=	167	;
						10'd491	:	dt	<=	201	;
						10'd492	:	dt	<=	202	;
						10'd493	:	dt	<=	210	;
						10'd494	:	dt	<=	200	;
						10'd495	:	dt	<=	185	;
						10'd496	:	dt	<=	165	;
						10'd497	:	dt	<=	134	;
						10'd498	:	dt	<=	88	;
						10'd499	:	dt	<=	134	;
						10'd500	:	dt	<=	221	;
						10'd501	:	dt	<=	207	;
						10'd502	:	dt	<=	208	;
						10'd503	:	dt	<=	207	;
						10'd504	:	dt	<=	216	;
						10'd505	:	dt	<=	216	;
						10'd506	:	dt	<=	217	;
						10'd507	:	dt	<=	217	;
						10'd508	:	dt	<=	217	;
						10'd509	:	dt	<=	217	;
						10'd510	:	dt	<=	217	;
						10'd511	:	dt	<=	195	;
						10'd512	:	dt	<=	199	;
						10'd513	:	dt	<=	195	;
						10'd514	:	dt	<=	159	;
						10'd515	:	dt	<=	132	;
						10'd516	:	dt	<=	126	;
						10'd517	:	dt	<=	129	;
						10'd518	:	dt	<=	176	;
						10'd519	:	dt	<=	207	;
						10'd520	:	dt	<=	211	;
						10'd521	:	dt	<=	210	;
						10'd522	:	dt	<=	192	;
						10'd523	:	dt	<=	173	;
						10'd524	:	dt	<=	155	;
						10'd525	:	dt	<=	118	;
						10'd526	:	dt	<=	80	;
						10'd527	:	dt	<=	183	;
						10'd528	:	dt	<=	218	;
						10'd529	:	dt	<=	209	;
						10'd530	:	dt	<=	209	;
						10'd531	:	dt	<=	208	;
						10'd532	:	dt	<=	217	;
						10'd533	:	dt	<=	217	;
						10'd534	:	dt	<=	218	;
						10'd535	:	dt	<=	218	;
						10'd536	:	dt	<=	218	;
						10'd537	:	dt	<=	218	;
						10'd538	:	dt	<=	220	;
						10'd539	:	dt	<=	195	;
						10'd540	:	dt	<=	193	;
						10'd541	:	dt	<=	196	;
						10'd542	:	dt	<=	169	;
						10'd543	:	dt	<=	139	;
						10'd544	:	dt	<=	128	;
						10'd545	:	dt	<=	134	;
						10'd546	:	dt	<=	183	;
						10'd547	:	dt	<=	212	;
						10'd548	:	dt	<=	211	;
						10'd549	:	dt	<=	202	;
						10'd550	:	dt	<=	184	;
						10'd551	:	dt	<=	164	;
						10'd552	:	dt	<=	147	;
						10'd553	:	dt	<=	100	;
						10'd554	:	dt	<=	101	;
						10'd555	:	dt	<=	217	;
						10'd556	:	dt	<=	211	;
						10'd557	:	dt	<=	211	;
						10'd558	:	dt	<=	210	;
						10'd559	:	dt	<=	209	;
						10'd560	:	dt	<=	217	;
						10'd561	:	dt	<=	217	;
						10'd562	:	dt	<=	218	;
						10'd563	:	dt	<=	219	;
						10'd564	:	dt	<=	218	;
						10'd565	:	dt	<=	218	;
						10'd566	:	dt	<=	221	;
						10'd567	:	dt	<=	199	;
						10'd568	:	dt	<=	180	;
						10'd569	:	dt	<=	187	;
						10'd570	:	dt	<=	169	;
						10'd571	:	dt	<=	142	;
						10'd572	:	dt	<=	129	;
						10'd573	:	dt	<=	140	;
						10'd574	:	dt	<=	192	;
						10'd575	:	dt	<=	209	;
						10'd576	:	dt	<=	200	;
						10'd577	:	dt	<=	193	;
						10'd578	:	dt	<=	174	;
						10'd579	:	dt	<=	150	;
						10'd580	:	dt	<=	134	;
						10'd581	:	dt	<=	85	;
						10'd582	:	dt	<=	150	;
						10'd583	:	dt	<=	224	;
						10'd584	:	dt	<=	209	;
						10'd585	:	dt	<=	212	;
						10'd586	:	dt	<=	210	;
						10'd587	:	dt	<=	210	;
						10'd588	:	dt	<=	217	;
						10'd589	:	dt	<=	217	;
						10'd590	:	dt	<=	217	;
						10'd591	:	dt	<=	218	;
						10'd592	:	dt	<=	218	;
						10'd593	:	dt	<=	218	;
						10'd594	:	dt	<=	221	;
						10'd595	:	dt	<=	212	;
						10'd596	:	dt	<=	177	;
						10'd597	:	dt	<=	187	;
						10'd598	:	dt	<=	175	;
						10'd599	:	dt	<=	145	;
						10'd600	:	dt	<=	139	;
						10'd601	:	dt	<=	145	;
						10'd602	:	dt	<=	196	;
						10'd603	:	dt	<=	200	;
						10'd604	:	dt	<=	191	;
						10'd605	:	dt	<=	182	;
						10'd606	:	dt	<=	161	;
						10'd607	:	dt	<=	137	;
						10'd608	:	dt	<=	113	;
						10'd609	:	dt	<=	85	;
						10'd610	:	dt	<=	201	;
						10'd611	:	dt	<=	219	;
						10'd612	:	dt	<=	213	;
						10'd613	:	dt	<=	212	;
						10'd614	:	dt	<=	211	;
						10'd615	:	dt	<=	211	;
						10'd616	:	dt	<=	216	;
						10'd617	:	dt	<=	216	;
						10'd618	:	dt	<=	217	;
						10'd619	:	dt	<=	218	;
						10'd620	:	dt	<=	217	;
						10'd621	:	dt	<=	217	;
						10'd622	:	dt	<=	217	;
						10'd623	:	dt	<=	220	;
						10'd624	:	dt	<=	189	;
						10'd625	:	dt	<=	185	;
						10'd626	:	dt	<=	180	;
						10'd627	:	dt	<=	159	;
						10'd628	:	dt	<=	157	;
						10'd629	:	dt	<=	142	;
						10'd630	:	dt	<=	192	;
						10'd631	:	dt	<=	191	;
						10'd632	:	dt	<=	188	;
						10'd633	:	dt	<=	168	;
						10'd634	:	dt	<=	146	;
						10'd635	:	dt	<=	127	;
						10'd636	:	dt	<=	87	;
						10'd637	:	dt	<=	125	;
						10'd638	:	dt	<=	225	;
						10'd639	:	dt	<=	212	;
						10'd640	:	dt	<=	214	;
						10'd641	:	dt	<=	212	;
						10'd642	:	dt	<=	210	;
						10'd643	:	dt	<=	210	;
						10'd644	:	dt	<=	216	;
						10'd645	:	dt	<=	216	;
						10'd646	:	dt	<=	217	;
						10'd647	:	dt	<=	218	;
						10'd648	:	dt	<=	217	;
						10'd649	:	dt	<=	217	;
						10'd650	:	dt	<=	217	;
						10'd651	:	dt	<=	222	;
						10'd652	:	dt	<=	204	;
						10'd653	:	dt	<=	181	;
						10'd654	:	dt	<=	181	;
						10'd655	:	dt	<=	171	;
						10'd656	:	dt	<=	157	;
						10'd657	:	dt	<=	133	;
						10'd658	:	dt	<=	174	;
						10'd659	:	dt	<=	182	;
						10'd660	:	dt	<=	179	;
						10'd661	:	dt	<=	156	;
						10'd662	:	dt	<=	128	;
						10'd663	:	dt	<=	106	;
						10'd664	:	dt	<=	79	;
						10'd665	:	dt	<=	194	;
						10'd666	:	dt	<=	218	;
						10'd667	:	dt	<=	211	;
						10'd668	:	dt	<=	211	;
						10'd669	:	dt	<=	211	;
						10'd670	:	dt	<=	210	;
						10'd671	:	dt	<=	210	;
						10'd672	:	dt	<=	217	;
						10'd673	:	dt	<=	216	;
						10'd674	:	dt	<=	218	;
						10'd675	:	dt	<=	218	;
						10'd676	:	dt	<=	218	;
						10'd677	:	dt	<=	218	;
						10'd678	:	dt	<=	218	;
						10'd679	:	dt	<=	221	;
						10'd680	:	dt	<=	211	;
						10'd681	:	dt	<=	186	;
						10'd682	:	dt	<=	178	;
						10'd683	:	dt	<=	165	;
						10'd684	:	dt	<=	151	;
						10'd685	:	dt	<=	135	;
						10'd686	:	dt	<=	156	;
						10'd687	:	dt	<=	164	;
						10'd688	:	dt	<=	153	;
						10'd689	:	dt	<=	130	;
						10'd690	:	dt	<=	107	;
						10'd691	:	dt	<=	73	;
						10'd692	:	dt	<=	141	;
						10'd693	:	dt	<=	226	;
						10'd694	:	dt	<=	212	;
						10'd695	:	dt	<=	214	;
						10'd696	:	dt	<=	213	;
						10'd697	:	dt	<=	212	;
						10'd698	:	dt	<=	211	;
						10'd699	:	dt	<=	210	;
						10'd700	:	dt	<=	217	;
						10'd701	:	dt	<=	218	;
						10'd702	:	dt	<=	218	;
						10'd703	:	dt	<=	218	;
						10'd704	:	dt	<=	218	;
						10'd705	:	dt	<=	218	;
						10'd706	:	dt	<=	219	;
						10'd707	:	dt	<=	221	;
						10'd708	:	dt	<=	213	;
						10'd709	:	dt	<=	193	;
						10'd710	:	dt	<=	181	;
						10'd711	:	dt	<=	163	;
						10'd712	:	dt	<=	148	;
						10'd713	:	dt	<=	137	;
						10'd714	:	dt	<=	145	;
						10'd715	:	dt	<=	154	;
						10'd716	:	dt	<=	133	;
						10'd717	:	dt	<=	108	;
						10'd718	:	dt	<=	84	;
						10'd719	:	dt	<=	89	;
						10'd720	:	dt	<=	213	;
						10'd721	:	dt	<=	218	;
						10'd722	:	dt	<=	216	;
						10'd723	:	dt	<=	215	;
						10'd724	:	dt	<=	213	;
						10'd725	:	dt	<=	212	;
						10'd726	:	dt	<=	211	;
						10'd727	:	dt	<=	210	;
						10'd728	:	dt	<=	217	;
						10'd729	:	dt	<=	219	;
						10'd730	:	dt	<=	219	;
						10'd731	:	dt	<=	219	;
						10'd732	:	dt	<=	218	;
						10'd733	:	dt	<=	218	;
						10'd734	:	dt	<=	220	;
						10'd735	:	dt	<=	222	;
						10'd736	:	dt	<=	203	;
						10'd737	:	dt	<=	194	;
						10'd738	:	dt	<=	182	;
						10'd739	:	dt	<=	167	;
						10'd740	:	dt	<=	155	;
						10'd741	:	dt	<=	148	;
						10'd742	:	dt	<=	143	;
						10'd743	:	dt	<=	149	;
						10'd744	:	dt	<=	136	;
						10'd745	:	dt	<=	106	;
						10'd746	:	dt	<=	72	;
						10'd747	:	dt	<=	150	;
						10'd748	:	dt	<=	229	;
						10'd749	:	dt	<=	214	;
						10'd750	:	dt	<=	217	;
						10'd751	:	dt	<=	215	;
						10'd752	:	dt	<=	213	;
						10'd753	:	dt	<=	212	;
						10'd754	:	dt	<=	211	;
						10'd755	:	dt	<=	212	;
						10'd756	:	dt	<=	217	;
						10'd757	:	dt	<=	217	;
						10'd758	:	dt	<=	218	;
						10'd759	:	dt	<=	218	;
						10'd760	:	dt	<=	219	;
						10'd761	:	dt	<=	218	;
						10'd762	:	dt	<=	220	;
						10'd763	:	dt	<=	218	;
						10'd764	:	dt	<=	190	;
						10'd765	:	dt	<=	193	;
						10'd766	:	dt	<=	185	;
						10'd767	:	dt	<=	178	;
						10'd768	:	dt	<=	175	;
						10'd769	:	dt	<=	162	;
						10'd770	:	dt	<=	150	;
						10'd771	:	dt	<=	142	;
						10'd772	:	dt	<=	128	;
						10'd773	:	dt	<=	97	;
						10'd774	:	dt	<=	81	;
						10'd775	:	dt	<=	192	;
						10'd776	:	dt	<=	223	;
						10'd777	:	dt	<=	216	;
						10'd778	:	dt	<=	216	;
						10'd779	:	dt	<=	215	;
						10'd780	:	dt	<=	214	;
						10'd781	:	dt	<=	213	;
						10'd782	:	dt	<=	212	;
						10'd783	:	dt	<=	204	;
					endcase
				end
				5'd5	:	begin
					case (cnt)
						10'd0	:	dt	<=	126	;
						10'd1	:	dt	<=	128	;
						10'd2	:	dt	<=	131	;
						10'd3	:	dt	<=	132	;
						10'd4	:	dt	<=	133	;
						10'd5	:	dt	<=	134	;
						10'd6	:	dt	<=	135	;
						10'd7	:	dt	<=	135	;
						10'd8	:	dt	<=	136	;
						10'd9	:	dt	<=	138	;
						10'd10	:	dt	<=	137	;
						10'd11	:	dt	<=	137	;
						10'd12	:	dt	<=	138	;
						10'd13	:	dt	<=	138	;
						10'd14	:	dt	<=	139	;
						10'd15	:	dt	<=	137	;
						10'd16	:	dt	<=	142	;
						10'd17	:	dt	<=	140	;
						10'd18	:	dt	<=	138	;
						10'd19	:	dt	<=	139	;
						10'd20	:	dt	<=	137	;
						10'd21	:	dt	<=	137	;
						10'd22	:	dt	<=	136	;
						10'd23	:	dt	<=	135	;
						10'd24	:	dt	<=	134	;
						10'd25	:	dt	<=	133	;
						10'd26	:	dt	<=	134	;
						10'd27	:	dt	<=	132	;
						10'd28	:	dt	<=	129	;
						10'd29	:	dt	<=	132	;
						10'd30	:	dt	<=	134	;
						10'd31	:	dt	<=	135	;
						10'd32	:	dt	<=	135	;
						10'd33	:	dt	<=	137	;
						10'd34	:	dt	<=	139	;
						10'd35	:	dt	<=	139	;
						10'd36	:	dt	<=	139	;
						10'd37	:	dt	<=	140	;
						10'd38	:	dt	<=	141	;
						10'd39	:	dt	<=	141	;
						10'd40	:	dt	<=	142	;
						10'd41	:	dt	<=	143	;
						10'd42	:	dt	<=	142	;
						10'd43	:	dt	<=	142	;
						10'd44	:	dt	<=	116	;
						10'd45	:	dt	<=	138	;
						10'd46	:	dt	<=	141	;
						10'd47	:	dt	<=	140	;
						10'd48	:	dt	<=	141	;
						10'd49	:	dt	<=	140	;
						10'd50	:	dt	<=	139	;
						10'd51	:	dt	<=	138	;
						10'd52	:	dt	<=	137	;
						10'd53	:	dt	<=	136	;
						10'd54	:	dt	<=	136	;
						10'd55	:	dt	<=	134	;
						10'd56	:	dt	<=	133	;
						10'd57	:	dt	<=	135	;
						10'd58	:	dt	<=	138	;
						10'd59	:	dt	<=	139	;
						10'd60	:	dt	<=	139	;
						10'd61	:	dt	<=	141	;
						10'd62	:	dt	<=	142	;
						10'd63	:	dt	<=	143	;
						10'd64	:	dt	<=	142	;
						10'd65	:	dt	<=	143	;
						10'd66	:	dt	<=	145	;
						10'd67	:	dt	<=	145	;
						10'd68	:	dt	<=	143	;
						10'd69	:	dt	<=	145	;
						10'd70	:	dt	<=	145	;
						10'd71	:	dt	<=	158	;
						10'd72	:	dt	<=	94	;
						10'd73	:	dt	<=	118	;
						10'd74	:	dt	<=	151	;
						10'd75	:	dt	<=	143	;
						10'd76	:	dt	<=	144	;
						10'd77	:	dt	<=	144	;
						10'd78	:	dt	<=	142	;
						10'd79	:	dt	<=	141	;
						10'd80	:	dt	<=	141	;
						10'd81	:	dt	<=	140	;
						10'd82	:	dt	<=	139	;
						10'd83	:	dt	<=	138	;
						10'd84	:	dt	<=	137	;
						10'd85	:	dt	<=	139	;
						10'd86	:	dt	<=	142	;
						10'd87	:	dt	<=	142	;
						10'd88	:	dt	<=	142	;
						10'd89	:	dt	<=	144	;
						10'd90	:	dt	<=	146	;
						10'd91	:	dt	<=	146	;
						10'd92	:	dt	<=	146	;
						10'd93	:	dt	<=	147	;
						10'd94	:	dt	<=	147	;
						10'd95	:	dt	<=	147	;
						10'd96	:	dt	<=	148	;
						10'd97	:	dt	<=	117	;
						10'd98	:	dt	<=	128	;
						10'd99	:	dt	<=	168	;
						10'd100	:	dt	<=	101	;
						10'd101	:	dt	<=	98	;
						10'd102	:	dt	<=	157	;
						10'd103	:	dt	<=	146	;
						10'd104	:	dt	<=	147	;
						10'd105	:	dt	<=	146	;
						10'd106	:	dt	<=	146	;
						10'd107	:	dt	<=	145	;
						10'd108	:	dt	<=	144	;
						10'd109	:	dt	<=	143	;
						10'd110	:	dt	<=	142	;
						10'd111	:	dt	<=	141	;
						10'd112	:	dt	<=	140	;
						10'd113	:	dt	<=	142	;
						10'd114	:	dt	<=	145	;
						10'd115	:	dt	<=	146	;
						10'd116	:	dt	<=	147	;
						10'd117	:	dt	<=	148	;
						10'd118	:	dt	<=	149	;
						10'd119	:	dt	<=	149	;
						10'd120	:	dt	<=	149	;
						10'd121	:	dt	<=	151	;
						10'd122	:	dt	<=	151	;
						10'd123	:	dt	<=	149	;
						10'd124	:	dt	<=	161	;
						10'd125	:	dt	<=	114	;
						10'd126	:	dt	<=	99	;
						10'd127	:	dt	<=	174	;
						10'd128	:	dt	<=	99	;
						10'd129	:	dt	<=	84	;
						10'd130	:	dt	<=	162	;
						10'd131	:	dt	<=	149	;
						10'd132	:	dt	<=	151	;
						10'd133	:	dt	<=	149	;
						10'd134	:	dt	<=	148	;
						10'd135	:	dt	<=	147	;
						10'd136	:	dt	<=	146	;
						10'd137	:	dt	<=	146	;
						10'd138	:	dt	<=	145	;
						10'd139	:	dt	<=	144	;
						10'd140	:	dt	<=	143	;
						10'd141	:	dt	<=	145	;
						10'd142	:	dt	<=	149	;
						10'd143	:	dt	<=	150	;
						10'd144	:	dt	<=	150	;
						10'd145	:	dt	<=	151	;
						10'd146	:	dt	<=	153	;
						10'd147	:	dt	<=	153	;
						10'd148	:	dt	<=	154	;
						10'd149	:	dt	<=	153	;
						10'd150	:	dt	<=	154	;
						10'd151	:	dt	<=	152	;
						10'd152	:	dt	<=	167	;
						10'd153	:	dt	<=	126	;
						10'd154	:	dt	<=	88	;
						10'd155	:	dt	<=	169	;
						10'd156	:	dt	<=	99	;
						10'd157	:	dt	<=	87	;
						10'd158	:	dt	<=	164	;
						10'd159	:	dt	<=	152	;
						10'd160	:	dt	<=	153	;
						10'd161	:	dt	<=	152	;
						10'd162	:	dt	<=	151	;
						10'd163	:	dt	<=	150	;
						10'd164	:	dt	<=	149	;
						10'd165	:	dt	<=	148	;
						10'd166	:	dt	<=	148	;
						10'd167	:	dt	<=	147	;
						10'd168	:	dt	<=	145	;
						10'd169	:	dt	<=	147	;
						10'd170	:	dt	<=	151	;
						10'd171	:	dt	<=	152	;
						10'd172	:	dt	<=	153	;
						10'd173	:	dt	<=	155	;
						10'd174	:	dt	<=	155	;
						10'd175	:	dt	<=	155	;
						10'd176	:	dt	<=	151	;
						10'd177	:	dt	<=	154	;
						10'd178	:	dt	<=	158	;
						10'd179	:	dt	<=	155	;
						10'd180	:	dt	<=	170	;
						10'd181	:	dt	<=	130	;
						10'd182	:	dt	<=	79	;
						10'd183	:	dt	<=	166	;
						10'd184	:	dt	<=	111	;
						10'd185	:	dt	<=	93	;
						10'd186	:	dt	<=	166	;
						10'd187	:	dt	<=	156	;
						10'd188	:	dt	<=	157	;
						10'd189	:	dt	<=	156	;
						10'd190	:	dt	<=	155	;
						10'd191	:	dt	<=	153	;
						10'd192	:	dt	<=	152	;
						10'd193	:	dt	<=	152	;
						10'd194	:	dt	<=	152	;
						10'd195	:	dt	<=	150	;
						10'd196	:	dt	<=	149	;
						10'd197	:	dt	<=	150	;
						10'd198	:	dt	<=	153	;
						10'd199	:	dt	<=	155	;
						10'd200	:	dt	<=	155	;
						10'd201	:	dt	<=	158	;
						10'd202	:	dt	<=	157	;
						10'd203	:	dt	<=	163	;
						10'd204	:	dt	<=	129	;
						10'd205	:	dt	<=	120	;
						10'd206	:	dt	<=	166	;
						10'd207	:	dt	<=	156	;
						10'd208	:	dt	<=	171	;
						10'd209	:	dt	<=	140	;
						10'd210	:	dt	<=	82	;
						10'd211	:	dt	<=	162	;
						10'd212	:	dt	<=	102	;
						10'd213	:	dt	<=	97	;
						10'd214	:	dt	<=	168	;
						10'd215	:	dt	<=	158	;
						10'd216	:	dt	<=	160	;
						10'd217	:	dt	<=	158	;
						10'd218	:	dt	<=	162	;
						10'd219	:	dt	<=	160	;
						10'd220	:	dt	<=	154	;
						10'd221	:	dt	<=	154	;
						10'd222	:	dt	<=	154	;
						10'd223	:	dt	<=	152	;
						10'd224	:	dt	<=	151	;
						10'd225	:	dt	<=	152	;
						10'd226	:	dt	<=	156	;
						10'd227	:	dt	<=	158	;
						10'd228	:	dt	<=	159	;
						10'd229	:	dt	<=	159	;
						10'd230	:	dt	<=	158	;
						10'd231	:	dt	<=	164	;
						10'd232	:	dt	<=	139	;
						10'd233	:	dt	<=	91	;
						10'd234	:	dt	<=	165	;
						10'd235	:	dt	<=	159	;
						10'd236	:	dt	<=	174	;
						10'd237	:	dt	<=	144	;
						10'd238	:	dt	<=	71	;
						10'd239	:	dt	<=	156	;
						10'd240	:	dt	<=	96	;
						10'd241	:	dt	<=	100	;
						10'd242	:	dt	<=	171	;
						10'd243	:	dt	<=	161	;
						10'd244	:	dt	<=	161	;
						10'd245	:	dt	<=	158	;
						10'd246	:	dt	<=	128	;
						10'd247	:	dt	<=	145	;
						10'd248	:	dt	<=	162	;
						10'd249	:	dt	<=	156	;
						10'd250	:	dt	<=	155	;
						10'd251	:	dt	<=	155	;
						10'd252	:	dt	<=	152	;
						10'd253	:	dt	<=	155	;
						10'd254	:	dt	<=	159	;
						10'd255	:	dt	<=	160	;
						10'd256	:	dt	<=	161	;
						10'd257	:	dt	<=	161	;
						10'd258	:	dt	<=	160	;
						10'd259	:	dt	<=	168	;
						10'd260	:	dt	<=	158	;
						10'd261	:	dt	<=	76	;
						10'd262	:	dt	<=	159	;
						10'd263	:	dt	<=	164	;
						10'd264	:	dt	<=	172	;
						10'd265	:	dt	<=	142	;
						10'd266	:	dt	<=	63	;
						10'd267	:	dt	<=	155	;
						10'd268	:	dt	<=	117	;
						10'd269	:	dt	<=	100	;
						10'd270	:	dt	<=	174	;
						10'd271	:	dt	<=	159	;
						10'd272	:	dt	<=	164	;
						10'd273	:	dt	<=	164	;
						10'd274	:	dt	<=	126	;
						10'd275	:	dt	<=	103	;
						10'd276	:	dt	<=	162	;
						10'd277	:	dt	<=	161	;
						10'd278	:	dt	<=	158	;
						10'd279	:	dt	<=	157	;
						10'd280	:	dt	<=	153	;
						10'd281	:	dt	<=	157	;
						10'd282	:	dt	<=	160	;
						10'd283	:	dt	<=	162	;
						10'd284	:	dt	<=	162	;
						10'd285	:	dt	<=	162	;
						10'd286	:	dt	<=	164	;
						10'd287	:	dt	<=	167	;
						10'd288	:	dt	<=	158	;
						10'd289	:	dt	<=	78	;
						10'd290	:	dt	<=	158	;
						10'd291	:	dt	<=	167	;
						10'd292	:	dt	<=	167	;
						10'd293	:	dt	<=	156	;
						10'd294	:	dt	<=	73	;
						10'd295	:	dt	<=	133	;
						10'd296	:	dt	<=	129	;
						10'd297	:	dt	<=	102	;
						10'd298	:	dt	<=	172	;
						10'd299	:	dt	<=	157	;
						10'd300	:	dt	<=	148	;
						10'd301	:	dt	<=	130	;
						10'd302	:	dt	<=	156	;
						10'd303	:	dt	<=	132	;
						10'd304	:	dt	<=	129	;
						10'd305	:	dt	<=	163	;
						10'd306	:	dt	<=	161	;
						10'd307	:	dt	<=	159	;
						10'd308	:	dt	<=	157	;
						10'd309	:	dt	<=	159	;
						10'd310	:	dt	<=	162	;
						10'd311	:	dt	<=	164	;
						10'd312	:	dt	<=	164	;
						10'd313	:	dt	<=	165	;
						10'd314	:	dt	<=	166	;
						10'd315	:	dt	<=	167	;
						10'd316	:	dt	<=	173	;
						10'd317	:	dt	<=	89	;
						10'd318	:	dt	<=	139	;
						10'd319	:	dt	<=	172	;
						10'd320	:	dt	<=	162	;
						10'd321	:	dt	<=	163	;
						10'd322	:	dt	<=	79	;
						10'd323	:	dt	<=	98	;
						10'd324	:	dt	<=	132	;
						10'd325	:	dt	<=	111	;
						10'd326	:	dt	<=	170	;
						10'd327	:	dt	<=	160	;
						10'd328	:	dt	<=	142	;
						10'd329	:	dt	<=	54	;
						10'd330	:	dt	<=	125	;
						10'd331	:	dt	<=	150	;
						10'd332	:	dt	<=	102	;
						10'd333	:	dt	<=	150	;
						10'd334	:	dt	<=	167	;
						10'd335	:	dt	<=	162	;
						10'd336	:	dt	<=	159	;
						10'd337	:	dt	<=	161	;
						10'd338	:	dt	<=	166	;
						10'd339	:	dt	<=	165	;
						10'd340	:	dt	<=	167	;
						10'd341	:	dt	<=	167	;
						10'd342	:	dt	<=	167	;
						10'd343	:	dt	<=	168	;
						10'd344	:	dt	<=	178	;
						10'd345	:	dt	<=	118	;
						10'd346	:	dt	<=	112	;
						10'd347	:	dt	<=	175	;
						10'd348	:	dt	<=	164	;
						10'd349	:	dt	<=	167	;
						10'd350	:	dt	<=	82	;
						10'd351	:	dt	<=	91	;
						10'd352	:	dt	<=	129	;
						10'd353	:	dt	<=	110	;
						10'd354	:	dt	<=	160	;
						10'd355	:	dt	<=	156	;
						10'd356	:	dt	<=	130	;
						10'd357	:	dt	<=	96	;
						10'd358	:	dt	<=	157	;
						10'd359	:	dt	<=	130	;
						10'd360	:	dt	<=	106	;
						10'd361	:	dt	<=	169	;
						10'd362	:	dt	<=	165	;
						10'd363	:	dt	<=	164	;
						10'd364	:	dt	<=	159	;
						10'd365	:	dt	<=	162	;
						10'd366	:	dt	<=	166	;
						10'd367	:	dt	<=	167	;
						10'd368	:	dt	<=	168	;
						10'd369	:	dt	<=	168	;
						10'd370	:	dt	<=	170	;
						10'd371	:	dt	<=	169	;
						10'd372	:	dt	<=	164	;
						10'd373	:	dt	<=	168	;
						10'd374	:	dt	<=	132	;
						10'd375	:	dt	<=	141	;
						10'd376	:	dt	<=	162	;
						10'd377	:	dt	<=	153	;
						10'd378	:	dt	<=	103	;
						10'd379	:	dt	<=	113	;
						10'd380	:	dt	<=	117	;
						10'd381	:	dt	<=	96	;
						10'd382	:	dt	<=	133	;
						10'd383	:	dt	<=	143	;
						10'd384	:	dt	<=	107	;
						10'd385	:	dt	<=	147	;
						10'd386	:	dt	<=	172	;
						10'd387	:	dt	<=	99	;
						10'd388	:	dt	<=	139	;
						10'd389	:	dt	<=	174	;
						10'd390	:	dt	<=	165	;
						10'd391	:	dt	<=	166	;
						10'd392	:	dt	<=	161	;
						10'd393	:	dt	<=	164	;
						10'd394	:	dt	<=	167	;
						10'd395	:	dt	<=	170	;
						10'd396	:	dt	<=	171	;
						10'd397	:	dt	<=	171	;
						10'd398	:	dt	<=	170	;
						10'd399	:	dt	<=	173	;
						10'd400	:	dt	<=	160	;
						10'd401	:	dt	<=	173	;
						10'd402	:	dt	<=	162	;
						10'd403	:	dt	<=	129	;
						10'd404	:	dt	<=	132	;
						10'd405	:	dt	<=	132	;
						10'd406	:	dt	<=	109	;
						10'd407	:	dt	<=	109	;
						10'd408	:	dt	<=	108	;
						10'd409	:	dt	<=	99	;
						10'd410	:	dt	<=	135	;
						10'd411	:	dt	<=	142	;
						10'd412	:	dt	<=	111	;
						10'd413	:	dt	<=	163	;
						10'd414	:	dt	<=	154	;
						10'd415	:	dt	<=	77	;
						10'd416	:	dt	<=	156	;
						10'd417	:	dt	<=	172	;
						10'd418	:	dt	<=	167	;
						10'd419	:	dt	<=	167	;
						10'd420	:	dt	<=	165	;
						10'd421	:	dt	<=	167	;
						10'd422	:	dt	<=	168	;
						10'd423	:	dt	<=	171	;
						10'd424	:	dt	<=	172	;
						10'd425	:	dt	<=	173	;
						10'd426	:	dt	<=	173	;
						10'd427	:	dt	<=	174	;
						10'd428	:	dt	<=	169	;
						10'd429	:	dt	<=	170	;
						10'd430	:	dt	<=	182	;
						10'd431	:	dt	<=	150	;
						10'd432	:	dt	<=	125	;
						10'd433	:	dt	<=	124	;
						10'd434	:	dt	<=	100	;
						10'd435	:	dt	<=	106	;
						10'd436	:	dt	<=	103	;
						10'd437	:	dt	<=	102	;
						10'd438	:	dt	<=	130	;
						10'd439	:	dt	<=	138	;
						10'd440	:	dt	<=	124	;
						10'd441	:	dt	<=	178	;
						10'd442	:	dt	<=	130	;
						10'd443	:	dt	<=	64	;
						10'd444	:	dt	<=	168	;
						10'd445	:	dt	<=	172	;
						10'd446	:	dt	<=	170	;
						10'd447	:	dt	<=	169	;
						10'd448	:	dt	<=	165	;
						10'd449	:	dt	<=	168	;
						10'd450	:	dt	<=	170	;
						10'd451	:	dt	<=	171	;
						10'd452	:	dt	<=	172	;
						10'd453	:	dt	<=	174	;
						10'd454	:	dt	<=	175	;
						10'd455	:	dt	<=	174	;
						10'd456	:	dt	<=	175	;
						10'd457	:	dt	<=	172	;
						10'd458	:	dt	<=	195	;
						10'd459	:	dt	<=	170	;
						10'd460	:	dt	<=	114	;
						10'd461	:	dt	<=	110	;
						10'd462	:	dt	<=	94	;
						10'd463	:	dt	<=	89	;
						10'd464	:	dt	<=	98	;
						10'd465	:	dt	<=	105	;
						10'd466	:	dt	<=	127	;
						10'd467	:	dt	<=	134	;
						10'd468	:	dt	<=	124	;
						10'd469	:	dt	<=	182	;
						10'd470	:	dt	<=	126	;
						10'd471	:	dt	<=	80	;
						10'd472	:	dt	<=	180	;
						10'd473	:	dt	<=	171	;
						10'd474	:	dt	<=	171	;
						10'd475	:	dt	<=	171	;
						10'd476	:	dt	<=	166	;
						10'd477	:	dt	<=	169	;
						10'd478	:	dt	<=	171	;
						10'd479	:	dt	<=	172	;
						10'd480	:	dt	<=	173	;
						10'd481	:	dt	<=	174	;
						10'd482	:	dt	<=	175	;
						10'd483	:	dt	<=	176	;
						10'd484	:	dt	<=	177	;
						10'd485	:	dt	<=	174	;
						10'd486	:	dt	<=	197	;
						10'd487	:	dt	<=	179	;
						10'd488	:	dt	<=	119	;
						10'd489	:	dt	<=	86	;
						10'd490	:	dt	<=	87	;
						10'd491	:	dt	<=	81	;
						10'd492	:	dt	<=	94	;
						10'd493	:	dt	<=	118	;
						10'd494	:	dt	<=	136	;
						10'd495	:	dt	<=	123	;
						10'd496	:	dt	<=	116	;
						10'd497	:	dt	<=	177	;
						10'd498	:	dt	<=	127	;
						10'd499	:	dt	<=	94	;
						10'd500	:	dt	<=	183	;
						10'd501	:	dt	<=	172	;
						10'd502	:	dt	<=	173	;
						10'd503	:	dt	<=	173	;
						10'd504	:	dt	<=	169	;
						10'd505	:	dt	<=	172	;
						10'd506	:	dt	<=	172	;
						10'd507	:	dt	<=	174	;
						10'd508	:	dt	<=	175	;
						10'd509	:	dt	<=	174	;
						10'd510	:	dt	<=	177	;
						10'd511	:	dt	<=	178	;
						10'd512	:	dt	<=	178	;
						10'd513	:	dt	<=	175	;
						10'd514	:	dt	<=	192	;
						10'd515	:	dt	<=	176	;
						10'd516	:	dt	<=	126	;
						10'd517	:	dt	<=	87	;
						10'd518	:	dt	<=	86	;
						10'd519	:	dt	<=	82	;
						10'd520	:	dt	<=	109	;
						10'd521	:	dt	<=	130	;
						10'd522	:	dt	<=	147	;
						10'd523	:	dt	<=	159	;
						10'd524	:	dt	<=	128	;
						10'd525	:	dt	<=	164	;
						10'd526	:	dt	<=	128	;
						10'd527	:	dt	<=	100	;
						10'd528	:	dt	<=	184	;
						10'd529	:	dt	<=	174	;
						10'd530	:	dt	<=	173	;
						10'd531	:	dt	<=	173	;
						10'd532	:	dt	<=	169	;
						10'd533	:	dt	<=	172	;
						10'd534	:	dt	<=	173	;
						10'd535	:	dt	<=	173	;
						10'd536	:	dt	<=	176	;
						10'd537	:	dt	<=	178	;
						10'd538	:	dt	<=	179	;
						10'd539	:	dt	<=	178	;
						10'd540	:	dt	<=	181	;
						10'd541	:	dt	<=	175	;
						10'd542	:	dt	<=	189	;
						10'd543	:	dt	<=	171	;
						10'd544	:	dt	<=	126	;
						10'd545	:	dt	<=	89	;
						10'd546	:	dt	<=	80	;
						10'd547	:	dt	<=	90	;
						10'd548	:	dt	<=	121	;
						10'd549	:	dt	<=	137	;
						10'd550	:	dt	<=	164	;
						10'd551	:	dt	<=	175	;
						10'd552	:	dt	<=	141	;
						10'd553	:	dt	<=	140	;
						10'd554	:	dt	<=	108	;
						10'd555	:	dt	<=	95	;
						10'd556	:	dt	<=	184	;
						10'd557	:	dt	<=	176	;
						10'd558	:	dt	<=	175	;
						10'd559	:	dt	<=	173	;
						10'd560	:	dt	<=	171	;
						10'd561	:	dt	<=	173	;
						10'd562	:	dt	<=	174	;
						10'd563	:	dt	<=	175	;
						10'd564	:	dt	<=	177	;
						10'd565	:	dt	<=	179	;
						10'd566	:	dt	<=	179	;
						10'd567	:	dt	<=	179	;
						10'd568	:	dt	<=	181	;
						10'd569	:	dt	<=	174	;
						10'd570	:	dt	<=	189	;
						10'd571	:	dt	<=	171	;
						10'd572	:	dt	<=	134	;
						10'd573	:	dt	<=	91	;
						10'd574	:	dt	<=	80	;
						10'd575	:	dt	<=	98	;
						10'd576	:	dt	<=	134	;
						10'd577	:	dt	<=	159	;
						10'd578	:	dt	<=	164	;
						10'd579	:	dt	<=	167	;
						10'd580	:	dt	<=	153	;
						10'd581	:	dt	<=	114	;
						10'd582	:	dt	<=	73	;
						10'd583	:	dt	<=	82	;
						10'd584	:	dt	<=	185	;
						10'd585	:	dt	<=	176	;
						10'd586	:	dt	<=	177	;
						10'd587	:	dt	<=	177	;
						10'd588	:	dt	<=	172	;
						10'd589	:	dt	<=	173	;
						10'd590	:	dt	<=	174	;
						10'd591	:	dt	<=	177	;
						10'd592	:	dt	<=	178	;
						10'd593	:	dt	<=	179	;
						10'd594	:	dt	<=	180	;
						10'd595	:	dt	<=	180	;
						10'd596	:	dt	<=	183	;
						10'd597	:	dt	<=	174	;
						10'd598	:	dt	<=	186	;
						10'd599	:	dt	<=	172	;
						10'd600	:	dt	<=	138	;
						10'd601	:	dt	<=	93	;
						10'd602	:	dt	<=	82	;
						10'd603	:	dt	<=	97	;
						10'd604	:	dt	<=	143	;
						10'd605	:	dt	<=	172	;
						10'd606	:	dt	<=	169	;
						10'd607	:	dt	<=	160	;
						10'd608	:	dt	<=	132	;
						10'd609	:	dt	<=	89	;
						10'd610	:	dt	<=	44	;
						10'd611	:	dt	<=	108	;
						10'd612	:	dt	<=	189	;
						10'd613	:	dt	<=	176	;
						10'd614	:	dt	<=	178	;
						10'd615	:	dt	<=	178	;
						10'd616	:	dt	<=	171	;
						10'd617	:	dt	<=	173	;
						10'd618	:	dt	<=	177	;
						10'd619	:	dt	<=	178	;
						10'd620	:	dt	<=	179	;
						10'd621	:	dt	<=	180	;
						10'd622	:	dt	<=	181	;
						10'd623	:	dt	<=	182	;
						10'd624	:	dt	<=	185	;
						10'd625	:	dt	<=	178	;
						10'd626	:	dt	<=	179	;
						10'd627	:	dt	<=	170	;
						10'd628	:	dt	<=	137	;
						10'd629	:	dt	<=	95	;
						10'd630	:	dt	<=	88	;
						10'd631	:	dt	<=	90	;
						10'd632	:	dt	<=	152	;
						10'd633	:	dt	<=	180	;
						10'd634	:	dt	<=	167	;
						10'd635	:	dt	<=	141	;
						10'd636	:	dt	<=	112	;
						10'd637	:	dt	<=	65	;
						10'd638	:	dt	<=	64	;
						10'd639	:	dt	<=	176	;
						10'd640	:	dt	<=	183	;
						10'd641	:	dt	<=	179	;
						10'd642	:	dt	<=	179	;
						10'd643	:	dt	<=	178	;
						10'd644	:	dt	<=	173	;
						10'd645	:	dt	<=	174	;
						10'd646	:	dt	<=	178	;
						10'd647	:	dt	<=	179	;
						10'd648	:	dt	<=	179	;
						10'd649	:	dt	<=	180	;
						10'd650	:	dt	<=	182	;
						10'd651	:	dt	<=	183	;
						10'd652	:	dt	<=	186	;
						10'd653	:	dt	<=	175	;
						10'd654	:	dt	<=	165	;
						10'd655	:	dt	<=	168	;
						10'd656	:	dt	<=	137	;
						10'd657	:	dt	<=	100	;
						10'd658	:	dt	<=	96	;
						10'd659	:	dt	<=	88	;
						10'd660	:	dt	<=	149	;
						10'd661	:	dt	<=	168	;
						10'd662	:	dt	<=	147	;
						10'd663	:	dt	<=	122	;
						10'd664	:	dt	<=	92	;
						10'd665	:	dt	<=	50	;
						10'd666	:	dt	<=	144	;
						10'd667	:	dt	<=	193	;
						10'd668	:	dt	<=	181	;
						10'd669	:	dt	<=	181	;
						10'd670	:	dt	<=	180	;
						10'd671	:	dt	<=	179	;
						10'd672	:	dt	<=	173	;
						10'd673	:	dt	<=	174	;
						10'd674	:	dt	<=	177	;
						10'd675	:	dt	<=	179	;
						10'd676	:	dt	<=	180	;
						10'd677	:	dt	<=	180	;
						10'd678	:	dt	<=	183	;
						10'd679	:	dt	<=	182	;
						10'd680	:	dt	<=	187	;
						10'd681	:	dt	<=	177	;
						10'd682	:	dt	<=	158	;
						10'd683	:	dt	<=	161	;
						10'd684	:	dt	<=	130	;
						10'd685	:	dt	<=	111	;
						10'd686	:	dt	<=	101	;
						10'd687	:	dt	<=	91	;
						10'd688	:	dt	<=	136	;
						10'd689	:	dt	<=	150	;
						10'd690	:	dt	<=	135	;
						10'd691	:	dt	<=	112	;
						10'd692	:	dt	<=	62	;
						10'd693	:	dt	<=	87	;
						10'd694	:	dt	<=	192	;
						10'd695	:	dt	<=	183	;
						10'd696	:	dt	<=	185	;
						10'd697	:	dt	<=	183	;
						10'd698	:	dt	<=	181	;
						10'd699	:	dt	<=	180	;
						10'd700	:	dt	<=	173	;
						10'd701	:	dt	<=	174	;
						10'd702	:	dt	<=	177	;
						10'd703	:	dt	<=	178	;
						10'd704	:	dt	<=	179	;
						10'd705	:	dt	<=	179	;
						10'd706	:	dt	<=	181	;
						10'd707	:	dt	<=	182	;
						10'd708	:	dt	<=	184	;
						10'd709	:	dt	<=	179	;
						10'd710	:	dt	<=	156	;
						10'd711	:	dt	<=	151	;
						10'd712	:	dt	<=	124	;
						10'd713	:	dt	<=	116	;
						10'd714	:	dt	<=	96	;
						10'd715	:	dt	<=	88	;
						10'd716	:	dt	<=	128	;
						10'd717	:	dt	<=	138	;
						10'd718	:	dt	<=	126	;
						10'd719	:	dt	<=	81	;
						10'd720	:	dt	<=	49	;
						10'd721	:	dt	<=	164	;
						10'd722	:	dt	<=	190	;
						10'd723	:	dt	<=	184	;
						10'd724	:	dt	<=	185	;
						10'd725	:	dt	<=	184	;
						10'd726	:	dt	<=	182	;
						10'd727	:	dt	<=	181	;
						10'd728	:	dt	<=	172	;
						10'd729	:	dt	<=	174	;
						10'd730	:	dt	<=	177	;
						10'd731	:	dt	<=	178	;
						10'd732	:	dt	<=	178	;
						10'd733	:	dt	<=	178	;
						10'd734	:	dt	<=	180	;
						10'd735	:	dt	<=	182	;
						10'd736	:	dt	<=	184	;
						10'd737	:	dt	<=	177	;
						10'd738	:	dt	<=	160	;
						10'd739	:	dt	<=	154	;
						10'd740	:	dt	<=	128	;
						10'd741	:	dt	<=	114	;
						10'd742	:	dt	<=	97	;
						10'd743	:	dt	<=	78	;
						10'd744	:	dt	<=	114	;
						10'd745	:	dt	<=	112	;
						10'd746	:	dt	<=	89	;
						10'd747	:	dt	<=	48	;
						10'd748	:	dt	<=	133	;
						10'd749	:	dt	<=	194	;
						10'd750	:	dt	<=	182	;
						10'd751	:	dt	<=	185	;
						10'd752	:	dt	<=	184	;
						10'd753	:	dt	<=	184	;
						10'd754	:	dt	<=	182	;
						10'd755	:	dt	<=	181	;
						10'd756	:	dt	<=	172	;
						10'd757	:	dt	<=	174	;
						10'd758	:	dt	<=	177	;
						10'd759	:	dt	<=	178	;
						10'd760	:	dt	<=	178	;
						10'd761	:	dt	<=	179	;
						10'd762	:	dt	<=	181	;
						10'd763	:	dt	<=	183	;
						10'd764	:	dt	<=	187	;
						10'd765	:	dt	<=	175	;
						10'd766	:	dt	<=	165	;
						10'd767	:	dt	<=	154	;
						10'd768	:	dt	<=	118	;
						10'd769	:	dt	<=	107	;
						10'd770	:	dt	<=	100	;
						10'd771	:	dt	<=	75	;
						10'd772	:	dt	<=	96	;
						10'd773	:	dt	<=	83	;
						10'd774	:	dt	<=	47	;
						10'd775	:	dt	<=	104	;
						10'd776	:	dt	<=	194	;
						10'd777	:	dt	<=	183	;
						10'd778	:	dt	<=	186	;
						10'd779	:	dt	<=	184	;
						10'd780	:	dt	<=	184	;
						10'd781	:	dt	<=	184	;
						10'd782	:	dt	<=	182	;
						10'd783	:	dt	<=	180	;
					endcase
				end
				5'd14	:	begin
					case (cnt)
						10'd0	:	dt	<=	177	;
						10'd1	:	dt	<=	177	;
						10'd2	:	dt	<=	177	;
						10'd3	:	dt	<=	177	;
						10'd4	:	dt	<=	177	;
						10'd5	:	dt	<=	178	;
						10'd6	:	dt	<=	179	;
						10'd7	:	dt	<=	179	;
						10'd8	:	dt	<=	178	;
						10'd9	:	dt	<=	179	;
						10'd10	:	dt	<=	179	;
						10'd11	:	dt	<=	178	;
						10'd12	:	dt	<=	179	;
						10'd13	:	dt	<=	178	;
						10'd14	:	dt	<=	179	;
						10'd15	:	dt	<=	179	;
						10'd16	:	dt	<=	179	;
						10'd17	:	dt	<=	179	;
						10'd18	:	dt	<=	178	;
						10'd19	:	dt	<=	178	;
						10'd20	:	dt	<=	179	;
						10'd21	:	dt	<=	178	;
						10'd22	:	dt	<=	177	;
						10'd23	:	dt	<=	178	;
						10'd24	:	dt	<=	177	;
						10'd25	:	dt	<=	177	;
						10'd26	:	dt	<=	179	;
						10'd27	:	dt	<=	143	;
						10'd28	:	dt	<=	180	;
						10'd29	:	dt	<=	180	;
						10'd30	:	dt	<=	180	;
						10'd31	:	dt	<=	180	;
						10'd32	:	dt	<=	180	;
						10'd33	:	dt	<=	180	;
						10'd34	:	dt	<=	181	;
						10'd35	:	dt	<=	182	;
						10'd36	:	dt	<=	183	;
						10'd37	:	dt	<=	182	;
						10'd38	:	dt	<=	183	;
						10'd39	:	dt	<=	182	;
						10'd40	:	dt	<=	181	;
						10'd41	:	dt	<=	181	;
						10'd42	:	dt	<=	181	;
						10'd43	:	dt	<=	181	;
						10'd44	:	dt	<=	182	;
						10'd45	:	dt	<=	183	;
						10'd46	:	dt	<=	181	;
						10'd47	:	dt	<=	181	;
						10'd48	:	dt	<=	181	;
						10'd49	:	dt	<=	180	;
						10'd50	:	dt	<=	179	;
						10'd51	:	dt	<=	180	;
						10'd52	:	dt	<=	179	;
						10'd53	:	dt	<=	177	;
						10'd54	:	dt	<=	182	;
						10'd55	:	dt	<=	127	;
						10'd56	:	dt	<=	182	;
						10'd57	:	dt	<=	182	;
						10'd58	:	dt	<=	182	;
						10'd59	:	dt	<=	181	;
						10'd60	:	dt	<=	183	;
						10'd61	:	dt	<=	183	;
						10'd62	:	dt	<=	183	;
						10'd63	:	dt	<=	184	;
						10'd64	:	dt	<=	183	;
						10'd65	:	dt	<=	183	;
						10'd66	:	dt	<=	182	;
						10'd67	:	dt	<=	183	;
						10'd68	:	dt	<=	183	;
						10'd69	:	dt	<=	184	;
						10'd70	:	dt	<=	182	;
						10'd71	:	dt	<=	186	;
						10'd72	:	dt	<=	187	;
						10'd73	:	dt	<=	183	;
						10'd74	:	dt	<=	184	;
						10'd75	:	dt	<=	184	;
						10'd76	:	dt	<=	184	;
						10'd77	:	dt	<=	182	;
						10'd78	:	dt	<=	181	;
						10'd79	:	dt	<=	181	;
						10'd80	:	dt	<=	180	;
						10'd81	:	dt	<=	181	;
						10'd82	:	dt	<=	182	;
						10'd83	:	dt	<=	157	;
						10'd84	:	dt	<=	185	;
						10'd85	:	dt	<=	184	;
						10'd86	:	dt	<=	184	;
						10'd87	:	dt	<=	186	;
						10'd88	:	dt	<=	186	;
						10'd89	:	dt	<=	186	;
						10'd90	:	dt	<=	185	;
						10'd91	:	dt	<=	185	;
						10'd92	:	dt	<=	188	;
						10'd93	:	dt	<=	193	;
						10'd94	:	dt	<=	183	;
						10'd95	:	dt	<=	173	;
						10'd96	:	dt	<=	186	;
						10'd97	:	dt	<=	185	;
						10'd98	:	dt	<=	172	;
						10'd99	:	dt	<=	169	;
						10'd100	:	dt	<=	182	;
						10'd101	:	dt	<=	188	;
						10'd102	:	dt	<=	188	;
						10'd103	:	dt	<=	186	;
						10'd104	:	dt	<=	186	;
						10'd105	:	dt	<=	186	;
						10'd106	:	dt	<=	185	;
						10'd107	:	dt	<=	185	;
						10'd108	:	dt	<=	183	;
						10'd109	:	dt	<=	183	;
						10'd110	:	dt	<=	183	;
						10'd111	:	dt	<=	174	;
						10'd112	:	dt	<=	188	;
						10'd113	:	dt	<=	188	;
						10'd114	:	dt	<=	188	;
						10'd115	:	dt	<=	190	;
						10'd116	:	dt	<=	189	;
						10'd117	:	dt	<=	188	;
						10'd118	:	dt	<=	186	;
						10'd119	:	dt	<=	197	;
						10'd120	:	dt	<=	211	;
						10'd121	:	dt	<=	178	;
						10'd122	:	dt	<=	173	;
						10'd123	:	dt	<=	171	;
						10'd124	:	dt	<=	174	;
						10'd125	:	dt	<=	162	;
						10'd126	:	dt	<=	134	;
						10'd127	:	dt	<=	149	;
						10'd128	:	dt	<=	166	;
						10'd129	:	dt	<=	171	;
						10'd130	:	dt	<=	176	;
						10'd131	:	dt	<=	192	;
						10'd132	:	dt	<=	188	;
						10'd133	:	dt	<=	190	;
						10'd134	:	dt	<=	190	;
						10'd135	:	dt	<=	188	;
						10'd136	:	dt	<=	186	;
						10'd137	:	dt	<=	185	;
						10'd138	:	dt	<=	186	;
						10'd139	:	dt	<=	182	;
						10'd140	:	dt	<=	191	;
						10'd141	:	dt	<=	191	;
						10'd142	:	dt	<=	190	;
						10'd143	:	dt	<=	193	;
						10'd144	:	dt	<=	190	;
						10'd145	:	dt	<=	197	;
						10'd146	:	dt	<=	209	;
						10'd147	:	dt	<=	205	;
						10'd148	:	dt	<=	188	;
						10'd149	:	dt	<=	122	;
						10'd150	:	dt	<=	99	;
						10'd151	:	dt	<=	122	;
						10'd152	:	dt	<=	134	;
						10'd153	:	dt	<=	132	;
						10'd154	:	dt	<=	93	;
						10'd155	:	dt	<=	89	;
						10'd156	:	dt	<=	149	;
						10'd157	:	dt	<=	133	;
						10'd158	:	dt	<=	111	;
						10'd159	:	dt	<=	194	;
						10'd160	:	dt	<=	191	;
						10'd161	:	dt	<=	192	;
						10'd162	:	dt	<=	192	;
						10'd163	:	dt	<=	190	;
						10'd164	:	dt	<=	188	;
						10'd165	:	dt	<=	188	;
						10'd166	:	dt	<=	188	;
						10'd167	:	dt	<=	186	;
						10'd168	:	dt	<=	193	;
						10'd169	:	dt	<=	193	;
						10'd170	:	dt	<=	193	;
						10'd171	:	dt	<=	195	;
						10'd172	:	dt	<=	188	;
						10'd173	:	dt	<=	211	;
						10'd174	:	dt	<=	220	;
						10'd175	:	dt	<=	146	;
						10'd176	:	dt	<=	113	;
						10'd177	:	dt	<=	90	;
						10'd178	:	dt	<=	54	;
						10'd179	:	dt	<=	68	;
						10'd180	:	dt	<=	86	;
						10'd181	:	dt	<=	93	;
						10'd182	:	dt	<=	74	;
						10'd183	:	dt	<=	68	;
						10'd184	:	dt	<=	100	;
						10'd185	:	dt	<=	103	;
						10'd186	:	dt	<=	73	;
						10'd187	:	dt	<=	172	;
						10'd188	:	dt	<=	202	;
						10'd189	:	dt	<=	194	;
						10'd190	:	dt	<=	188	;
						10'd191	:	dt	<=	192	;
						10'd192	:	dt	<=	191	;
						10'd193	:	dt	<=	190	;
						10'd194	:	dt	<=	190	;
						10'd195	:	dt	<=	190	;
						10'd196	:	dt	<=	195	;
						10'd197	:	dt	<=	194	;
						10'd198	:	dt	<=	194	;
						10'd199	:	dt	<=	197	;
						10'd200	:	dt	<=	188	;
						10'd201	:	dt	<=	220	;
						10'd202	:	dt	<=	213	;
						10'd203	:	dt	<=	136	;
						10'd204	:	dt	<=	71	;
						10'd205	:	dt	<=	61	;
						10'd206	:	dt	<=	55	;
						10'd207	:	dt	<=	50	;
						10'd208	:	dt	<=	57	;
						10'd209	:	dt	<=	64	;
						10'd210	:	dt	<=	67	;
						10'd211	:	dt	<=	61	;
						10'd212	:	dt	<=	71	;
						10'd213	:	dt	<=	80	;
						10'd214	:	dt	<=	94	;
						10'd215	:	dt	<=	107	;
						10'd216	:	dt	<=	172	;
						10'd217	:	dt	<=	170	;
						10'd218	:	dt	<=	142	;
						10'd219	:	dt	<=	155	;
						10'd220	:	dt	<=	195	;
						10'd221	:	dt	<=	190	;
						10'd222	:	dt	<=	192	;
						10'd223	:	dt	<=	192	;
						10'd224	:	dt	<=	197	;
						10'd225	:	dt	<=	196	;
						10'd226	:	dt	<=	197	;
						10'd227	:	dt	<=	199	;
						10'd228	:	dt	<=	190	;
						10'd229	:	dt	<=	226	;
						10'd230	:	dt	<=	208	;
						10'd231	:	dt	<=	151	;
						10'd232	:	dt	<=	90	;
						10'd233	:	dt	<=	65	;
						10'd234	:	dt	<=	62	;
						10'd235	:	dt	<=	57	;
						10'd236	:	dt	<=	56	;
						10'd237	:	dt	<=	55	;
						10'd238	:	dt	<=	64	;
						10'd239	:	dt	<=	61	;
						10'd240	:	dt	<=	62	;
						10'd241	:	dt	<=	97	;
						10'd242	:	dt	<=	142	;
						10'd243	:	dt	<=	108	;
						10'd244	:	dt	<=	86	;
						10'd245	:	dt	<=	164	;
						10'd246	:	dt	<=	138	;
						10'd247	:	dt	<=	140	;
						10'd248	:	dt	<=	201	;
						10'd249	:	dt	<=	193	;
						10'd250	:	dt	<=	195	;
						10'd251	:	dt	<=	193	;
						10'd252	:	dt	<=	200	;
						10'd253	:	dt	<=	198	;
						10'd254	:	dt	<=	200	;
						10'd255	:	dt	<=	199	;
						10'd256	:	dt	<=	192	;
						10'd257	:	dt	<=	227	;
						10'd258	:	dt	<=	194	;
						10'd259	:	dt	<=	128	;
						10'd260	:	dt	<=	71	;
						10'd261	:	dt	<=	55	;
						10'd262	:	dt	<=	61	;
						10'd263	:	dt	<=	70	;
						10'd264	:	dt	<=	67	;
						10'd265	:	dt	<=	55	;
						10'd266	:	dt	<=	65	;
						10'd267	:	dt	<=	69	;
						10'd268	:	dt	<=	64	;
						10'd269	:	dt	<=	78	;
						10'd270	:	dt	<=	97	;
						10'd271	:	dt	<=	71	;
						10'd272	:	dt	<=	136	;
						10'd273	:	dt	<=	185	;
						10'd274	:	dt	<=	110	;
						10'd275	:	dt	<=	164	;
						10'd276	:	dt	<=	205	;
						10'd277	:	dt	<=	196	;
						10'd278	:	dt	<=	197	;
						10'd279	:	dt	<=	196	;
						10'd280	:	dt	<=	200	;
						10'd281	:	dt	<=	199	;
						10'd282	:	dt	<=	201	;
						10'd283	:	dt	<=	199	;
						10'd284	:	dt	<=	203	;
						10'd285	:	dt	<=	228	;
						10'd286	:	dt	<=	191	;
						10'd287	:	dt	<=	148	;
						10'd288	:	dt	<=	104	;
						10'd289	:	dt	<=	68	;
						10'd290	:	dt	<=	55	;
						10'd291	:	dt	<=	67	;
						10'd292	:	dt	<=	59	;
						10'd293	:	dt	<=	71	;
						10'd294	:	dt	<=	63	;
						10'd295	:	dt	<=	86	;
						10'd296	:	dt	<=	138	;
						10'd297	:	dt	<=	173	;
						10'd298	:	dt	<=	151	;
						10'd299	:	dt	<=	120	;
						10'd300	:	dt	<=	185	;
						10'd301	:	dt	<=	172	;
						10'd302	:	dt	<=	100	;
						10'd303	:	dt	<=	175	;
						10'd304	:	dt	<=	206	;
						10'd305	:	dt	<=	198	;
						10'd306	:	dt	<=	198	;
						10'd307	:	dt	<=	198	;
						10'd308	:	dt	<=	202	;
						10'd309	:	dt	<=	202	;
						10'd310	:	dt	<=	203	;
						10'd311	:	dt	<=	200	;
						10'd312	:	dt	<=	211	;
						10'd313	:	dt	<=	231	;
						10'd314	:	dt	<=	198	;
						10'd315	:	dt	<=	162	;
						10'd316	:	dt	<=	127	;
						10'd317	:	dt	<=	93	;
						10'd318	:	dt	<=	78	;
						10'd319	:	dt	<=	59	;
						10'd320	:	dt	<=	62	;
						10'd321	:	dt	<=	94	;
						10'd322	:	dt	<=	72	;
						10'd323	:	dt	<=	135	;
						10'd324	:	dt	<=	220	;
						10'd325	:	dt	<=	205	;
						10'd326	:	dt	<=	213	;
						10'd327	:	dt	<=	191	;
						10'd328	:	dt	<=	189	;
						10'd329	:	dt	<=	170	;
						10'd330	:	dt	<=	98	;
						10'd331	:	dt	<=	169	;
						10'd332	:	dt	<=	208	;
						10'd333	:	dt	<=	199	;
						10'd334	:	dt	<=	200	;
						10'd335	:	dt	<=	200	;
						10'd336	:	dt	<=	205	;
						10'd337	:	dt	<=	205	;
						10'd338	:	dt	<=	206	;
						10'd339	:	dt	<=	200	;
						10'd340	:	dt	<=	218	;
						10'd341	:	dt	<=	237	;
						10'd342	:	dt	<=	207	;
						10'd343	:	dt	<=	167	;
						10'd344	:	dt	<=	115	;
						10'd345	:	dt	<=	90	;
						10'd346	:	dt	<=	82	;
						10'd347	:	dt	<=	76	;
						10'd348	:	dt	<=	76	;
						10'd349	:	dt	<=	80	;
						10'd350	:	dt	<=	74	;
						10'd351	:	dt	<=	175	;
						10'd352	:	dt	<=	211	;
						10'd353	:	dt	<=	202	;
						10'd354	:	dt	<=	204	;
						10'd355	:	dt	<=	177	;
						10'd356	:	dt	<=	185	;
						10'd357	:	dt	<=	161	;
						10'd358	:	dt	<=	99	;
						10'd359	:	dt	<=	158	;
						10'd360	:	dt	<=	212	;
						10'd361	:	dt	<=	200	;
						10'd362	:	dt	<=	201	;
						10'd363	:	dt	<=	201	;
						10'd364	:	dt	<=	205	;
						10'd365	:	dt	<=	206	;
						10'd366	:	dt	<=	207	;
						10'd367	:	dt	<=	201	;
						10'd368	:	dt	<=	221	;
						10'd369	:	dt	<=	243	;
						10'd370	:	dt	<=	213	;
						10'd371	:	dt	<=	168	;
						10'd372	:	dt	<=	108	;
						10'd373	:	dt	<=	83	;
						10'd374	:	dt	<=	77	;
						10'd375	:	dt	<=	74	;
						10'd376	:	dt	<=	91	;
						10'd377	:	dt	<=	76	;
						10'd378	:	dt	<=	97	;
						10'd379	:	dt	<=	212	;
						10'd380	:	dt	<=	205	;
						10'd381	:	dt	<=	208	;
						10'd382	:	dt	<=	197	;
						10'd383	:	dt	<=	183	;
						10'd384	:	dt	<=	187	;
						10'd385	:	dt	<=	156	;
						10'd386	:	dt	<=	98	;
						10'd387	:	dt	<=	135	;
						10'd388	:	dt	<=	216	;
						10'd389	:	dt	<=	202	;
						10'd390	:	dt	<=	202	;
						10'd391	:	dt	<=	202	;
						10'd392	:	dt	<=	206	;
						10'd393	:	dt	<=	207	;
						10'd394	:	dt	<=	207	;
						10'd395	:	dt	<=	204	;
						10'd396	:	dt	<=	222	;
						10'd397	:	dt	<=	242	;
						10'd398	:	dt	<=	215	;
						10'd399	:	dt	<=	181	;
						10'd400	:	dt	<=	131	;
						10'd401	:	dt	<=	89	;
						10'd402	:	dt	<=	69	;
						10'd403	:	dt	<=	70	;
						10'd404	:	dt	<=	88	;
						10'd405	:	dt	<=	74	;
						10'd406	:	dt	<=	129	;
						10'd407	:	dt	<=	222	;
						10'd408	:	dt	<=	203	;
						10'd409	:	dt	<=	209	;
						10'd410	:	dt	<=	187	;
						10'd411	:	dt	<=	199	;
						10'd412	:	dt	<=	191	;
						10'd413	:	dt	<=	149	;
						10'd414	:	dt	<=	86	;
						10'd415	:	dt	<=	163	;
						10'd416	:	dt	<=	215	;
						10'd417	:	dt	<=	203	;
						10'd418	:	dt	<=	205	;
						10'd419	:	dt	<=	204	;
						10'd420	:	dt	<=	206	;
						10'd421	:	dt	<=	207	;
						10'd422	:	dt	<=	210	;
						10'd423	:	dt	<=	203	;
						10'd424	:	dt	<=	220	;
						10'd425	:	dt	<=	245	;
						10'd426	:	dt	<=	218	;
						10'd427	:	dt	<=	183	;
						10'd428	:	dt	<=	144	;
						10'd429	:	dt	<=	101	;
						10'd430	:	dt	<=	70	;
						10'd431	:	dt	<=	68	;
						10'd432	:	dt	<=	81	;
						10'd433	:	dt	<=	63	;
						10'd434	:	dt	<=	147	;
						10'd435	:	dt	<=	212	;
						10'd436	:	dt	<=	211	;
						10'd437	:	dt	<=	200	;
						10'd438	:	dt	<=	176	;
						10'd439	:	dt	<=	201	;
						10'd440	:	dt	<=	192	;
						10'd441	:	dt	<=	125	;
						10'd442	:	dt	<=	110	;
						10'd443	:	dt	<=	214	;
						10'd444	:	dt	<=	208	;
						10'd445	:	dt	<=	207	;
						10'd446	:	dt	<=	207	;
						10'd447	:	dt	<=	206	;
						10'd448	:	dt	<=	209	;
						10'd449	:	dt	<=	210	;
						10'd450	:	dt	<=	213	;
						10'd451	:	dt	<=	201	;
						10'd452	:	dt	<=	214	;
						10'd453	:	dt	<=	244	;
						10'd454	:	dt	<=	220	;
						10'd455	:	dt	<=	191	;
						10'd456	:	dt	<=	154	;
						10'd457	:	dt	<=	106	;
						10'd458	:	dt	<=	77	;
						10'd459	:	dt	<=	72	;
						10'd460	:	dt	<=	69	;
						10'd461	:	dt	<=	67	;
						10'd462	:	dt	<=	109	;
						10'd463	:	dt	<=	130	;
						10'd464	:	dt	<=	171	;
						10'd465	:	dt	<=	169	;
						10'd466	:	dt	<=	178	;
						10'd467	:	dt	<=	191	;
						10'd468	:	dt	<=	173	;
						10'd469	:	dt	<=	102	;
						10'd470	:	dt	<=	171	;
						10'd471	:	dt	<=	219	;
						10'd472	:	dt	<=	207	;
						10'd473	:	dt	<=	210	;
						10'd474	:	dt	<=	207	;
						10'd475	:	dt	<=	207	;
						10'd476	:	dt	<=	211	;
						10'd477	:	dt	<=	211	;
						10'd478	:	dt	<=	213	;
						10'd479	:	dt	<=	202	;
						10'd480	:	dt	<=	214	;
						10'd481	:	dt	<=	243	;
						10'd482	:	dt	<=	221	;
						10'd483	:	dt	<=	193	;
						10'd484	:	dt	<=	162	;
						10'd485	:	dt	<=	121	;
						10'd486	:	dt	<=	86	;
						10'd487	:	dt	<=	57	;
						10'd488	:	dt	<=	72	;
						10'd489	:	dt	<=	84	;
						10'd490	:	dt	<=	100	;
						10'd491	:	dt	<=	128	;
						10'd492	:	dt	<=	146	;
						10'd493	:	dt	<=	156	;
						10'd494	:	dt	<=	173	;
						10'd495	:	dt	<=	177	;
						10'd496	:	dt	<=	139	;
						10'd497	:	dt	<=	113	;
						10'd498	:	dt	<=	211	;
						10'd499	:	dt	<=	211	;
						10'd500	:	dt	<=	212	;
						10'd501	:	dt	<=	213	;
						10'd502	:	dt	<=	211	;
						10'd503	:	dt	<=	209	;
						10'd504	:	dt	<=	211	;
						10'd505	:	dt	<=	211	;
						10'd506	:	dt	<=	214	;
						10'd507	:	dt	<=	204	;
						10'd508	:	dt	<=	215	;
						10'd509	:	dt	<=	242	;
						10'd510	:	dt	<=	226	;
						10'd511	:	dt	<=	196	;
						10'd512	:	dt	<=	167	;
						10'd513	:	dt	<=	133	;
						10'd514	:	dt	<=	100	;
						10'd515	:	dt	<=	59	;
						10'd516	:	dt	<=	77	;
						10'd517	:	dt	<=	90	;
						10'd518	:	dt	<=	120	;
						10'd519	:	dt	<=	148	;
						10'd520	:	dt	<=	159	;
						10'd521	:	dt	<=	155	;
						10'd522	:	dt	<=	150	;
						10'd523	:	dt	<=	150	;
						10'd524	:	dt	<=	106	;
						10'd525	:	dt	<=	158	;
						10'd526	:	dt	<=	222	;
						10'd527	:	dt	<=	212	;
						10'd528	:	dt	<=	214	;
						10'd529	:	dt	<=	214	;
						10'd530	:	dt	<=	212	;
						10'd531	:	dt	<=	210	;
						10'd532	:	dt	<=	213	;
						10'd533	:	dt	<=	212	;
						10'd534	:	dt	<=	215	;
						10'd535	:	dt	<=	203	;
						10'd536	:	dt	<=	213	;
						10'd537	:	dt	<=	241	;
						10'd538	:	dt	<=	227	;
						10'd539	:	dt	<=	201	;
						10'd540	:	dt	<=	172	;
						10'd541	:	dt	<=	138	;
						10'd542	:	dt	<=	108	;
						10'd543	:	dt	<=	72	;
						10'd544	:	dt	<=	76	;
						10'd545	:	dt	<=	104	;
						10'd546	:	dt	<=	139	;
						10'd547	:	dt	<=	161	;
						10'd548	:	dt	<=	164	;
						10'd549	:	dt	<=	144	;
						10'd550	:	dt	<=	130	;
						10'd551	:	dt	<=	114	;
						10'd552	:	dt	<=	94	;
						10'd553	:	dt	<=	204	;
						10'd554	:	dt	<=	217	;
						10'd555	:	dt	<=	215	;
						10'd556	:	dt	<=	214	;
						10'd557	:	dt	<=	214	;
						10'd558	:	dt	<=	213	;
						10'd559	:	dt	<=	213	;
						10'd560	:	dt	<=	214	;
						10'd561	:	dt	<=	212	;
						10'd562	:	dt	<=	216	;
						10'd563	:	dt	<=	203	;
						10'd564	:	dt	<=	206	;
						10'd565	:	dt	<=	240	;
						10'd566	:	dt	<=	225	;
						10'd567	:	dt	<=	205	;
						10'd568	:	dt	<=	175	;
						10'd569	:	dt	<=	143	;
						10'd570	:	dt	<=	111	;
						10'd571	:	dt	<=	87	;
						10'd572	:	dt	<=	75	;
						10'd573	:	dt	<=	103	;
						10'd574	:	dt	<=	142	;
						10'd575	:	dt	<=	161	;
						10'd576	:	dt	<=	161	;
						10'd577	:	dt	<=	141	;
						10'd578	:	dt	<=	112	;
						10'd579	:	dt	<=	93	;
						10'd580	:	dt	<=	121	;
						10'd581	:	dt	<=	225	;
						10'd582	:	dt	<=	212	;
						10'd583	:	dt	<=	214	;
						10'd584	:	dt	<=	214	;
						10'd585	:	dt	<=	215	;
						10'd586	:	dt	<=	216	;
						10'd587	:	dt	<=	215	;
						10'd588	:	dt	<=	215	;
						10'd589	:	dt	<=	213	;
						10'd590	:	dt	<=	217	;
						10'd591	:	dt	<=	206	;
						10'd592	:	dt	<=	204	;
						10'd593	:	dt	<=	236	;
						10'd594	:	dt	<=	225	;
						10'd595	:	dt	<=	208	;
						10'd596	:	dt	<=	179	;
						10'd597	:	dt	<=	150	;
						10'd598	:	dt	<=	115	;
						10'd599	:	dt	<=	97	;
						10'd600	:	dt	<=	77	;
						10'd601	:	dt	<=	94	;
						10'd602	:	dt	<=	139	;
						10'd603	:	dt	<=	160	;
						10'd604	:	dt	<=	155	;
						10'd605	:	dt	<=	127	;
						10'd606	:	dt	<=	102	;
						10'd607	:	dt	<=	95	;
						10'd608	:	dt	<=	192	;
						10'd609	:	dt	<=	221	;
						10'd610	:	dt	<=	216	;
						10'd611	:	dt	<=	216	;
						10'd612	:	dt	<=	215	;
						10'd613	:	dt	<=	215	;
						10'd614	:	dt	<=	215	;
						10'd615	:	dt	<=	214	;
						10'd616	:	dt	<=	217	;
						10'd617	:	dt	<=	217	;
						10'd618	:	dt	<=	217	;
						10'd619	:	dt	<=	205	;
						10'd620	:	dt	<=	208	;
						10'd621	:	dt	<=	233	;
						10'd622	:	dt	<=	225	;
						10'd623	:	dt	<=	209	;
						10'd624	:	dt	<=	183	;
						10'd625	:	dt	<=	157	;
						10'd626	:	dt	<=	123	;
						10'd627	:	dt	<=	106	;
						10'd628	:	dt	<=	89	;
						10'd629	:	dt	<=	90	;
						10'd630	:	dt	<=	145	;
						10'd631	:	dt	<=	157	;
						10'd632	:	dt	<=	145	;
						10'd633	:	dt	<=	118	;
						10'd634	:	dt	<=	85	;
						10'd635	:	dt	<=	144	;
						10'd636	:	dt	<=	231	;
						10'd637	:	dt	<=	216	;
						10'd638	:	dt	<=	218	;
						10'd639	:	dt	<=	217	;
						10'd640	:	dt	<=	216	;
						10'd641	:	dt	<=	216	;
						10'd642	:	dt	<=	216	;
						10'd643	:	dt	<=	215	;
						10'd644	:	dt	<=	219	;
						10'd645	:	dt	<=	218	;
						10'd646	:	dt	<=	220	;
						10'd647	:	dt	<=	203	;
						10'd648	:	dt	<=	212	;
						10'd649	:	dt	<=	238	;
						10'd650	:	dt	<=	224	;
						10'd651	:	dt	<=	207	;
						10'd652	:	dt	<=	189	;
						10'd653	:	dt	<=	164	;
						10'd654	:	dt	<=	123	;
						10'd655	:	dt	<=	111	;
						10'd656	:	dt	<=	104	;
						10'd657	:	dt	<=	85	;
						10'd658	:	dt	<=	142	;
						10'd659	:	dt	<=	142	;
						10'd660	:	dt	<=	128	;
						10'd661	:	dt	<=	109	;
						10'd662	:	dt	<=	80	;
						10'd663	:	dt	<=	191	;
						10'd664	:	dt	<=	227	;
						10'd665	:	dt	<=	218	;
						10'd666	:	dt	<=	219	;
						10'd667	:	dt	<=	219	;
						10'd668	:	dt	<=	217	;
						10'd669	:	dt	<=	217	;
						10'd670	:	dt	<=	218	;
						10'd671	:	dt	<=	217	;
						10'd672	:	dt	<=	219	;
						10'd673	:	dt	<=	219	;
						10'd674	:	dt	<=	224	;
						10'd675	:	dt	<=	204	;
						10'd676	:	dt	<=	218	;
						10'd677	:	dt	<=	241	;
						10'd678	:	dt	<=	221	;
						10'd679	:	dt	<=	207	;
						10'd680	:	dt	<=	195	;
						10'd681	:	dt	<=	168	;
						10'd682	:	dt	<=	127	;
						10'd683	:	dt	<=	112	;
						10'd684	:	dt	<=	107	;
						10'd685	:	dt	<=	88	;
						10'd686	:	dt	<=	122	;
						10'd687	:	dt	<=	128	;
						10'd688	:	dt	<=	121	;
						10'd689	:	dt	<=	96	;
						10'd690	:	dt	<=	104	;
						10'd691	:	dt	<=	224	;
						10'd692	:	dt	<=	222	;
						10'd693	:	dt	<=	220	;
						10'd694	:	dt	<=	219	;
						10'd695	:	dt	<=	219	;
						10'd696	:	dt	<=	219	;
						10'd697	:	dt	<=	218	;
						10'd698	:	dt	<=	218	;
						10'd699	:	dt	<=	217	;
						10'd700	:	dt	<=	220	;
						10'd701	:	dt	<=	219	;
						10'd702	:	dt	<=	222	;
						10'd703	:	dt	<=	205	;
						10'd704	:	dt	<=	231	;
						10'd705	:	dt	<=	237	;
						10'd706	:	dt	<=	224	;
						10'd707	:	dt	<=	219	;
						10'd708	:	dt	<=	196	;
						10'd709	:	dt	<=	169	;
						10'd710	:	dt	<=	128	;
						10'd711	:	dt	<=	111	;
						10'd712	:	dt	<=	103	;
						10'd713	:	dt	<=	92	;
						10'd714	:	dt	<=	108	;
						10'd715	:	dt	<=	115	;
						10'd716	:	dt	<=	112	;
						10'd717	:	dt	<=	80	;
						10'd718	:	dt	<=	166	;
						10'd719	:	dt	<=	233	;
						10'd720	:	dt	<=	222	;
						10'd721	:	dt	<=	222	;
						10'd722	:	dt	<=	221	;
						10'd723	:	dt	<=	220	;
						10'd724	:	dt	<=	219	;
						10'd725	:	dt	<=	218	;
						10'd726	:	dt	<=	218	;
						10'd727	:	dt	<=	218	;
						10'd728	:	dt	<=	220	;
						10'd729	:	dt	<=	220	;
						10'd730	:	dt	<=	216	;
						10'd731	:	dt	<=	204	;
						10'd732	:	dt	<=	239	;
						10'd733	:	dt	<=	238	;
						10'd734	:	dt	<=	227	;
						10'd735	:	dt	<=	214	;
						10'd736	:	dt	<=	187	;
						10'd737	:	dt	<=	154	;
						10'd738	:	dt	<=	121	;
						10'd739	:	dt	<=	106	;
						10'd740	:	dt	<=	99	;
						10'd741	:	dt	<=	94	;
						10'd742	:	dt	<=	101	;
						10'd743	:	dt	<=	103	;
						10'd744	:	dt	<=	92	;
						10'd745	:	dt	<=	118	;
						10'd746	:	dt	<=	225	;
						10'd747	:	dt	<=	225	;
						10'd748	:	dt	<=	223	;
						10'd749	:	dt	<=	223	;
						10'd750	:	dt	<=	222	;
						10'd751	:	dt	<=	220	;
						10'd752	:	dt	<=	220	;
						10'd753	:	dt	<=	220	;
						10'd754	:	dt	<=	219	;
						10'd755	:	dt	<=	219	;
						10'd756	:	dt	<=	221	;
						10'd757	:	dt	<=	222	;
						10'd758	:	dt	<=	209	;
						10'd759	:	dt	<=	205	;
						10'd760	:	dt	<=	234	;
						10'd761	:	dt	<=	235	;
						10'd762	:	dt	<=	224	;
						10'd763	:	dt	<=	199	;
						10'd764	:	dt	<=	167	;
						10'd765	:	dt	<=	137	;
						10'd766	:	dt	<=	113	;
						10'd767	:	dt	<=	100	;
						10'd768	:	dt	<=	94	;
						10'd769	:	dt	<=	98	;
						10'd770	:	dt	<=	100	;
						10'd771	:	dt	<=	100	;
						10'd772	:	dt	<=	94	;
						10'd773	:	dt	<=	198	;
						10'd774	:	dt	<=	232	;
						10'd775	:	dt	<=	223	;
						10'd776	:	dt	<=	224	;
						10'd777	:	dt	<=	224	;
						10'd778	:	dt	<=	223	;
						10'd779	:	dt	<=	221	;
						10'd780	:	dt	<=	221	;
						10'd781	:	dt	<=	221	;
						10'd782	:	dt	<=	220	;
						10'd783	:	dt	<=	219	;
					endcase
				end
			endcase
		end
	end

	assign	q_data = dt;
	
endmodule
