`include "global.sv"
`include "timescale.sv"
module wieght_conv2_rom(
	input			clk,
	input			rstn,
	input	[11:0]	aa,
	input			cena,
	output reg		[`WDP_WEIGHT*`OUTPUT_NUM_CONV1*`OUTPUT_NUM_CONV2 -1:0]	qa
	);
	
	
	logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][`WDP_WEIGHT-1:0] weight	 = {
18'd7291,  18'd18863,  18'd12748,  18'd2984,  -18'd2274,  18'd14137,  
-18'd5319,  -18'd14541,  -18'd25492,  18'd6231,  18'd5735,  18'd8019,  
18'd1339,  -18'd9333,  -18'd11008,  -18'd4636,  18'd6547,  -18'd3472,  
18'd19144,  18'd30244,  18'd19099,  18'd14793,  -18'd1815,  -18'd3255,  
-18'd2923,  18'd6405,  -18'd7473,  -18'd2318,  -18'd6138,  -18'd3445,  
-18'd7322,  -18'd24200,  -18'd7184,  18'd4464,  18'd6645,  -18'd18787,  
18'd3950,  18'd9235,  18'd4222,  -18'd19995,  -18'd8736,  18'd6609,  
-18'd8043,  -18'd11289,  -18'd26406,  -18'd312,  18'd13920,  18'd10194,  
18'd175,  -18'd20428,  -18'd11734,  18'd6211,  18'd747,  -18'd5888,  
-18'd1022,  18'd5698,  18'd514,  -18'd7508,  -18'd3140,  -18'd6991,  
18'd1333,  18'd7413,  18'd18952,  -18'd1421,  18'd362,  -18'd1274,  
18'd122,  -18'd16809,  18'd2891,  -18'd25085,  -18'd6905,  -18'd18952,  
-18'd7888,  -18'd6738,  -18'd3012,  -18'd4069,  -18'd3829,  -18'd7127,  
-18'd13577,  -18'd15960,  -18'd3665,  18'd11654,  18'd1456,  -18'd6498,  
18'd15317,  18'd1750,  -18'd3341,  -18'd4889,  -18'd6237,  18'd17161,  
18'd15779,  18'd9079,  -18'd6929,  18'd112,  18'd10380,  -18'd6567,  

-18'd7030,  -18'd1718,  18'd13301,  18'd24607,  18'd2342,  18'd1260,  
18'd2914,  -18'd10157,  -18'd28550,  -18'd15118,  18'd9850,  -18'd11831,  
18'd5481,  -18'd3717,  -18'd29258,  -18'd16596,  18'd672,  18'd13711,  
-18'd4758,  18'd9129,  18'd20946,  -18'd10320,  18'd666,  -18'd10344,  
-18'd1788,  18'd1000,  -18'd3612,  -18'd1195,  18'd4566,  -18'd2157,  
18'd9392,  -18'd13022,  -18'd5544,  -18'd28757,  18'd10571,  -18'd16621,  
-18'd4897,  -18'd8688,  -18'd4815,  18'd15252,  18'd5156,  18'd25788,  
-18'd509,  -18'd10049,  -18'd42035,  -18'd18495,  18'd11129,  -18'd10014,  
18'd16444,  18'd8267,  -18'd7675,  18'd15100,  18'd479,  18'd6133,  
-18'd756,  18'd10442,  18'd13715,  18'd4278,  -18'd12287,  -18'd7752,  
18'd3662,  18'd7386,  18'd20758,  -18'd14136,  -18'd5612,  18'd10948,  
18'd638,  18'd30618,  18'd30513,  18'd14146,  -18'd7372,  18'd25967,  
-18'd6979,  18'd4233,  18'd1577,  -18'd5443,  -18'd6292,  -18'd3377,  
-18'd1564,  -18'd1671,  -18'd7353,  -18'd18401,  -18'd1014,  -18'd3556,  
18'd17449,  18'd14406,  18'd27030,  18'd6310,  -18'd6096,  18'd18660,  
18'd16110,  -18'd9154,  -18'd4910,  18'd36,  -18'd4321,  -18'd28394,  

-18'd19117,  -18'd683,  18'd6356,  18'd13936,  18'd6988,  18'd11051,  
18'd14824,  -18'd763,  -18'd743,  -18'd13432,  18'd3906,  -18'd27928,  
-18'd12796,  -18'd3196,  -18'd18293,  -18'd7989,  -18'd3757,  -18'd22199,  
-18'd12645,  -18'd33474,  -18'd75,  -18'd5556,  -18'd1931,  -18'd5161,  
18'd1596,  18'd6074,  18'd1892,  18'd4593,  -18'd2010,  -18'd971,  
18'd25570,  18'd663,  -18'd963,  -18'd7974,  18'd3386,  -18'd16593,  
-18'd1138,  -18'd40474,  -18'd28243,  -18'd8080,  -18'd304,  18'd2793,  
18'd3059,  -18'd12076,  -18'd31033,  -18'd14218,  18'd7342,  -18'd13043,  
18'd35286,  18'd22083,  18'd16582,  18'd715,  -18'd3654,  -18'd10874,  
-18'd24667,  -18'd16388,  18'd10980,  18'd21895,  18'd7393,  18'd19162,  
-18'd6997,  -18'd5051,  18'd21051,  18'd20798,  -18'd3884,  18'd47663,  
-18'd17246,  -18'd27008,  -18'd20871,  18'd5656,  18'd2482,  18'd23069,  
18'd529,  -18'd2907,  -18'd9397,  18'd57,  -18'd2088,  -18'd2416,  
18'd8605,  18'd18909,  18'd12731,  -18'd1934,  -18'd9438,  -18'd3514,  
18'd5317,  18'd17160,  18'd38164,  18'd15906,  18'd1470,  18'd24054,  
18'd4682,  -18'd5360,  18'd822,  -18'd17415,  18'd491,  -18'd37877,  

18'd10093,  18'd12195,  18'd8696,  -18'd7288,  18'd5022,  -18'd10687,  
18'd11298,  -18'd4494,  -18'd5999,  -18'd25731,  18'd4524,  -18'd22867,  
18'd7528,  -18'd19578,  -18'd8758,  -18'd8661,  18'd4495,  -18'd45787,  
-18'd37598,  -18'd48407,  -18'd16522,  -18'd5286,  18'd3673,  18'd1145,  
-18'd2580,  -18'd1880,  18'd1614,  -18'd752,  -18'd7019,  18'd1157,  
18'd36031,  18'd21461,  18'd31747,  -18'd14640,  -18'd12983,  -18'd28075,  
18'd5170,  18'd21972,  18'd17719,  -18'd9308,  -18'd5112,  18'd2324,  
18'd12352,  18'd7981,  -18'd16344,  -18'd38631,  -18'd2566,  -18'd19306,  
18'd16808,  18'd37598,  18'd19405,  -18'd4311,  -18'd12502,  18'd31381,  
18'd2075,  -18'd15913,  18'd15758,  18'd33760,  -18'd735,  -18'd28112,  
-18'd21820,  -18'd32029,  -18'd32924,  18'd45293,  18'd530,  18'd25984,  
18'd14289,  18'd16937,  18'd4007,  -18'd13790,  -18'd6581,  18'd11252,  
18'd3114,  -18'd6576,  -18'd8425,  -18'd8987,  -18'd2101,  -18'd1078,  
-18'd1249,  18'd11095,  18'd284,  18'd9504,  -18'd12146,  -18'd18263,  
-18'd5634,  -18'd808,  -18'd408,  18'd27270,  -18'd5812,  18'd32268,  
18'd1642,  -18'd9771,  -18'd3083,  -18'd18716,  -18'd9009,  -18'd47606,  

18'd419,  18'd23813,  18'd26240,  18'd5165,  -18'd7377,  18'd15768,  
-18'd2235,  18'd2075,  18'd10355,  -18'd15503,  -18'd3058,  -18'd14171,  
18'd26519,  -18'd2034,  18'd23787,  -18'd24343,  -18'd12371,  -18'd34104,  
-18'd20332,  -18'd30037,  -18'd37663,  -18'd54,  18'd18115,  18'd1670,  
-18'd6950,  -18'd6949,  -18'd324,  -18'd1521,  18'd1813,  -18'd5800,  
-18'd1935,  18'd6427,  18'd26570,  18'd17798,  -18'd15704,  18'd18899,  
-18'd1249,  -18'd1742,  18'd1269,  -18'd11215,  18'd952,  18'd15098,  
18'd15729,  -18'd683,  -18'd12181,  -18'd28537,  -18'd2798,  18'd5388,  
-18'd19904,  -18'd8101,  -18'd10660,  18'd1909,  -18'd9438,  18'd18088,  
18'd15831,  18'd34965,  18'd50591,  18'd22596,  18'd2956,  18'd23662,  
18'd3317,  18'd12309,  18'd12826,  -18'd8024,  -18'd716,  18'd11973,  
18'd13776,  18'd32622,  18'd19770,  18'd4459,  -18'd10133,  18'd19448,  
-18'd1323,  18'd363,  -18'd4883,  18'd211,  18'd2069,  18'd2593,  
-18'd19118,  18'd17896,  18'd25723,  18'd13049,  18'd3266,  -18'd8870,  
-18'd19383,  -18'd15237,  18'd11143,  18'd5696,  18'd177,  18'd40191,  
-18'd7566,  -18'd10676,  18'd23000,  18'd9899,  -18'd8478,  -18'd30025,  


18'd14381,  18'd29704,  18'd22626,  -18'd8389,  -18'd2711,  -18'd2496,  
-18'd10293,  -18'd7523,  -18'd26448,  18'd14849,  18'd15315,  18'd2752,  
-18'd5633,  -18'd12285,  -18'd14734,  18'd2744,  18'd7528,  -18'd5034,  
18'd18648,  18'd36800,  18'd32247,  18'd28874,  18'd289,  18'd24724,  
-18'd1331,  -18'd2665,  18'd1750,  18'd1047,  -18'd6912,  18'd3355,  
18'd3374,  -18'd8258,  -18'd573,  -18'd7697,  18'd7589,  -18'd25178,  
-18'd5715,  18'd11823,  18'd7551,  -18'd18540,  -18'd3159,  -18'd8199,  
-18'd8684,  18'd2817,  -18'd2729,  18'd16629,  18'd13610,  18'd5638,  
-18'd10927,  -18'd25355,  -18'd12298,  -18'd1031,  18'd5950,  18'd1511,  
-18'd23527,  -18'd14863,  18'd1852,  -18'd16973,  -18'd4469,  -18'd4466,  
18'd2425,  -18'd5493,  -18'd2329,  -18'd16013,  -18'd8278,  18'd16424,  
18'd3878,  -18'd9172,  -18'd7737,  -18'd24126,  -18'd1371,  -18'd6090,  
-18'd8209,  -18'd7662,  18'd4095,  -18'd7634,  -18'd4668,  -18'd4355,  
-18'd14540,  -18'd1221,  -18'd14887,  18'd21047,  -18'd407,  -18'd2520,  
-18'd1831,  -18'd21171,  -18'd18746,  -18'd1232,  -18'd3099,  18'd8690,  
18'd17086,  18'd15792,  -18'd12325,  18'd1691,  18'd10248,  -18'd4966,  

-18'd8326,  18'd13837,  18'd958,  18'd15472,  -18'd3687,  -18'd924,  
18'd5006,  18'd3313,  -18'd7529,  -18'd17629,  18'd10258,  -18'd15099,  
18'd4718,  -18'd16440,  -18'd659,  -18'd12467,  -18'd4105,  18'd4984,  
-18'd7931,  18'd21972,  18'd29319,  18'd23926,  -18'd7501,  18'd24535,  
18'd6850,  -18'd5081,  18'd4773,  -18'd5572,  -18'd262,  18'd1058,  
-18'd14703,  -18'd15548,  18'd8166,  -18'd1119,  -18'd1230,  -18'd445,  
-18'd19650,  -18'd36683,  -18'd15502,  -18'd224,  18'd2879,  18'd5768,  
18'd590,  -18'd23773,  -18'd31897,  -18'd10567,  18'd10362,  -18'd17026,  
18'd19133,  18'd9606,  -18'd4025,  18'd3166,  18'd8637,  -18'd439,  
-18'd5587,  18'd3197,  18'd6415,  18'd3577,  -18'd3302,  18'd15363,  
-18'd5155,  -18'd11663,  -18'd3674,  18'd19739,  -18'd5045,  18'd35223,  
-18'd6133,  18'd35246,  18'd19347,  18'd29259,  18'd2595,  18'd37675,  
-18'd6445,  -18'd4,  -18'd7701,  18'd4450,  -18'd1323,  -18'd3151,  
18'd18487,  -18'd1539,  18'd6685,  18'd5155,  -18'd2357,  -18'd25091,  
18'd14739,  18'd9685,  -18'd9926,  -18'd3939,  18'd5160,  18'd29385,  
18'd10743,  18'd16845,  -18'd936,  18'd994,  -18'd100,  -18'd7993,  

-18'd19344,  -18'd2483,  -18'd19809,  18'd15406,  -18'd277,  18'd12765,  
18'd12892,  18'd10749,  18'd8869,  -18'd30212,  -18'd973,  -18'd40315,  
18'd4044,  18'd605,  -18'd637,  -18'd19740,  -18'd4553,  -18'd18386,  
-18'd22280,  -18'd17311,  18'd9163,  18'd14694,  -18'd5956,  -18'd3133,  
-18'd4755,  18'd1726,  -18'd4527,  -18'd30,  18'd5396,  -18'd6874,  
18'd12177,  -18'd2063,  -18'd10857,  18'd2987,  -18'd2950,  -18'd7672,  
-18'd451,  -18'd50868,  -18'd25599,  -18'd22074,  18'd846,  -18'd29397,  
18'd4417,  -18'd1158,  -18'd15122,  -18'd29588,  18'd8114,  -18'd14138,  
18'd28874,  18'd15231,  18'd16656,  18'd647,  18'd2430,  -18'd9695,  
-18'd13225,  -18'd7979,  -18'd3999,  18'd36382,  -18'd1233,  18'd23169,  
-18'd8563,  -18'd7600,  -18'd33538,  18'd1259,  18'd8186,  18'd34203,  
-18'd15037,  -18'd6913,  -18'd42007,  18'd11586,  18'd12060,  18'd17909,  
18'd2824,  18'd232,  18'd4489,  18'd2628,  -18'd3777,  18'd36,  
18'd9385,  18'd31130,  18'd16718,  18'd7807,  -18'd7700,  18'd6688,  
-18'd10662,  18'd14049,  18'd4337,  18'd13420,  -18'd760,  18'd44737,  
18'd14457,  -18'd2873,  18'd6886,  -18'd24189,  -18'd8898,  -18'd14875,  

18'd17436,  18'd4798,  -18'd8659,  -18'd11482,  -18'd5100,  -18'd15573,  
18'd19333,  18'd9306,  18'd4323,  -18'd22648,  -18'd881,  -18'd29253,  
18'd13580,  -18'd9464,  18'd2932,  -18'd4129,  -18'd949,  -18'd31503,  
-18'd35289,  -18'd22789,  18'd8096,  18'd19609,  18'd11118,  18'd5069,  
-18'd3869,  -18'd6808,  -18'd3250,  -18'd4618,  -18'd6046,  -18'd5128,  
18'd22512,  18'd40708,  18'd18808,  -18'd16551,  -18'd5558,  18'd17316,  
18'd15472,  18'd5429,  18'd22813,  -18'd39926,  -18'd8719,  -18'd33899,  
18'd13332,  -18'd1479,  -18'd746,  -18'd19772,  18'd1944,  -18'd22231,  
18'd9453,  18'd30405,  18'd12189,  18'd16446,  -18'd2906,  18'd23864,  
18'd8423,  18'd1085,  18'd36381,  -18'd9298,  -18'd324,  18'd6616,  
-18'd447,  -18'd23192,  -18'd44432,  18'd6168,  18'd3252,  18'd6559,  
18'd21678,  18'd20477,  18'd1359,  -18'd20624,  18'd476,  -18'd2924,  
-18'd2311,  18'd731,  18'd2620,  -18'd67,  18'd1687,  -18'd7036,  
18'd12569,  18'd24803,  18'd973,  18'd20542,  -18'd16255,  18'd2513,  
-18'd24836,  -18'd21005,  -18'd39434,  -18'd9087,  18'd8891,  18'd33653,  
-18'd2827,  18'd861,  18'd1063,  -18'd10548,  -18'd17629,  -18'd33358,  

18'd8252,  18'd30364,  18'd8720,  18'd1453,  -18'd429,  18'd15031,  
-18'd2007,  -18'd4555,  18'd12290,  -18'd7402,  -18'd7678,  -18'd31791,  
18'd19188,  -18'd2117,  18'd16690,  -18'd22025,  -18'd10171,  -18'd22829,  
-18'd24292,  -18'd20404,  -18'd6582,  18'd12417,  18'd18212,  18'd5555,  
18'd1771,  -18'd5706,  18'd223,  18'd2650,  18'd2204,  18'd1964,  
18'd533,  18'd14078,  18'd11021,  18'd16835,  -18'd15495,  18'd14773,  
18'd7911,  18'd4814,  18'd2421,  -18'd13928,  18'd2814,  -18'd8550,  
18'd19824,  -18'd957,  18'd2378,  -18'd12815,  -18'd2089,  -18'd5181,  
-18'd23907,  -18'd12777,  -18'd30571,  18'd1784,  -18'd1061,  18'd16652,  
-18'd16985,  18'd42241,  18'd33858,  18'd47777,  18'd1415,  18'd67441,  
18'd10807,  18'd27150,  18'd16718,  -18'd34244,  -18'd6591,  -18'd2369,  
18'd11559,  18'd35360,  18'd16806,  18'd3583,  -18'd5958,  18'd36138,  
-18'd1658,  18'd5278,  18'd4358,  -18'd6388,  -18'd4010,  18'd1908,  
-18'd2560,  18'd32390,  18'd23667,  18'd14733,  -18'd6896,  18'd14684,  
-18'd632,  -18'd20190,  -18'd38247,  -18'd10646,  18'd5609,  18'd34343,  
-18'd83,  18'd2831,  18'd23405,  -18'd1968,  -18'd12449,  18'd3705,  


18'd18578,  18'd20482,  18'd5843,  -18'd11039,  -18'd4823,  -18'd9074,  
18'd7330,  18'd5866,  18'd9207,  18'd1751,  18'd11204,  -18'd13187,  
-18'd8923,  -18'd10032,  -18'd12261,  -18'd2146,  18'd1658,  18'd8701,  
18'd6592,  18'd30119,  18'd3634,  18'd3404,  -18'd8354,  18'd17156,  
-18'd2828,  -18'd1090,  -18'd2802,  18'd3763,  18'd77,  -18'd2886,  
-18'd2516,  -18'd4747,  18'd16242,  18'd8869,  -18'd1881,  -18'd4311,  
-18'd4458,  -18'd3899,  -18'd1324,  -18'd26174,  -18'd5399,  -18'd11404,  
-18'd11963,  -18'd5583,  18'd7683,  18'd25394,  18'd8115,  18'd10353,  
-18'd1380,  -18'd6806,  -18'd4028,  18'd13827,  18'd2109,  -18'd4983,  
-18'd25779,  -18'd21551,  -18'd6026,  -18'd14948,  18'd859,  -18'd7201,  
-18'd9986,  -18'd19253,  18'd2197,  -18'd3068,  18'd6190,  18'd1994,  
18'd2808,  -18'd8098,  18'd4659,  -18'd459,  -18'd2123,  -18'd3641,  
-18'd5366,  -18'd7885,  18'd3172,  -18'd2141,  -18'd7356,  -18'd6006,  
18'd100,  18'd12704,  18'd12065,  18'd31050,  18'd2348,  -18'd944,  
-18'd23871,  -18'd27012,  -18'd29490,  -18'd5242,  18'd12270,  18'd6763,  
18'd15081,  18'd11792,  18'd2549,  18'd5914,  18'd397,  18'd2379,  

-18'd3970,  18'd18400,  18'd6903,  18'd7311,  -18'd4643,  18'd7092,  
18'd5081,  18'd6941,  18'd23770,  -18'd157,  18'd7429,  -18'd38644,  
18'd15397,  -18'd8364,  -18'd17225,  -18'd18545,  18'd5362,  18'd5412,  
18'd577,  18'd22075,  18'd14053,  18'd29689,  -18'd15589,  18'd23133,  
-18'd2685,  -18'd4463,  -18'd3216,  -18'd5659,  18'd5633,  -18'd2902,  
-18'd16423,  -18'd20603,  -18'd4877,  18'd21746,  18'd6435,  18'd7460,  
-18'd25656,  -18'd42398,  -18'd5661,  -18'd9751,  18'd3515,  -18'd87,  
18'd902,  -18'd10513,  -18'd12606,  18'd3036,  18'd10234,  -18'd30247,  
18'd8072,  18'd8176,  -18'd13042,  18'd7039,  -18'd1535,  -18'd16338,  
-18'd6727,  -18'd14238,  -18'd19918,  18'd5436,  18'd2568,  -18'd2420,  
-18'd24661,  -18'd22007,  -18'd11752,  18'd11763,  18'd8567,  18'd9888,  
-18'd3857,  18'd28491,  18'd5227,  18'd17912,  18'd3378,  18'd18484,  
-18'd6655,  -18'd8622,  -18'd5502,  -18'd7069,  18'd3847,  -18'd4453,  
18'd9971,  18'd11984,  18'd24913,  18'd25988,  -18'd7073,  -18'd4439,  
-18'd514,  -18'd3132,  -18'd21798,  -18'd25993,  18'd11693,  18'd544,  
18'd23469,  18'd21122,  -18'd149,  -18'd7843,  18'd3764,  18'd462,  

-18'd19909,  -18'd22698,  -18'd29333,  18'd14211,  -18'd1781,  -18'd1698,  
18'd8370,  18'd4044,  18'd14577,  -18'd10173,  -18'd6574,  -18'd30159,  
18'd17841,  18'd12053,  -18'd10467,  -18'd22081,  -18'd2063,  -18'd28147,  
-18'd20697,  -18'd13798,  18'd10452,  18'd17742,  -18'd5330,  -18'd290,  
18'd2405,  18'd2245,  18'd446,  -18'd5908,  -18'd6987,  18'd610,  
18'd14116,  18'd9461,  -18'd12592,  18'd21195,  18'd5043,  -18'd24570,  
-18'd2938,  -18'd31329,  -18'd14747,  -18'd15041,  18'd4388,  -18'd27233,  
18'd7342,  -18'd4398,  -18'd5683,  -18'd26499,  -18'd429,  -18'd30681,  
18'd29191,  18'd21750,  18'd9495,  18'd3233,  -18'd5253,  -18'd22931,  
18'd9070,  -18'd2236,  18'd11778,  -18'd112,  -18'd6846,  -18'd9869,  
18'd8580,  -18'd4739,  -18'd13240,  -18'd6530,  18'd8456,  -18'd3478,  
-18'd3262,  18'd6206,  -18'd21901,  18'd15367,  18'd5444,  -18'd6033,  
18'd3336,  -18'd6274,  -18'd4430,  -18'd3264,  -18'd3281,  18'd1386,  
18'd4729,  18'd17706,  18'd21123,  18'd39706,  -18'd10591,  18'd14949,  
-18'd6556,  -18'd5292,  18'd1926,  -18'd14010,  18'd1157,  18'd24602,  
18'd14188,  18'd13080,  18'd11406,  -18'd17652,  -18'd10517,  18'd16007,  

18'd8351,  -18'd3981,  -18'd96,  -18'd20504,  18'd6965,  -18'd25722,  
18'd13738,  18'd4969,  18'd6285,  18'd2826,  -18'd8935,  -18'd17185,  
18'd13726,  18'd10829,  18'd28555,  -18'd6336,  -18'd4376,  -18'd19474,  
-18'd29576,  -18'd19497,  -18'd7541,  18'd27012,  18'd5628,  18'd3466,  
18'd3572,  -18'd72,  -18'd5535,  18'd65,  18'd3431,  18'd5089,  
18'd14593,  18'd29080,  18'd4952,  -18'd18894,  -18'd3328,  -18'd3369,  
18'd21505,  18'd12818,  18'd2721,  -18'd33817,  -18'd4165,  -18'd20078,  
18'd4292,  -18'd15910,  18'd5331,  -18'd19999,  -18'd2323,  -18'd6045,  
-18'd15848,  18'd15624,  18'd5807,  18'd28623,  -18'd4388,  18'd19532,  
18'd16002,  18'd27988,  18'd35189,  -18'd10858,  18'd8404,  18'd29046,  
18'd17842,  -18'd5662,  -18'd4694,  -18'd11966,  -18'd5475,  -18'd39515,  
18'd28258,  18'd10539,  18'd21508,  -18'd33474,  18'd3847,  -18'd35494,  
-18'd929,  -18'd9,  18'd5342,  -18'd4328,  -18'd83,  -18'd2162,  
18'd6518,  18'd14329,  18'd9181,  18'd23578,  -18'd3410,  18'd7386,  
-18'd12552,  -18'd24584,  -18'd23856,  -18'd2075,  18'd7226,  -18'd3207,  
-18'd6288,  18'd1219,  -18'd8935,  18'd11208,  -18'd15867,  18'd12633,  

18'd13827,  18'd10184,  18'd8016,  -18'd2249,  18'd6428,  18'd1868,  
-18'd1723,  18'd5671,  18'd23221,  18'd13653,  -18'd11679,  -18'd13098,  
18'd3061,  -18'd878,  18'd15245,  18'd20649,  -18'd9198,  -18'd2007,  
-18'd20855,  -18'd18515,  18'd12559,  18'd23561,  18'd12223,  18'd15028,  
-18'd3849,  -18'd5068,  18'd2449,  -18'd2496,  -18'd3377,  18'd2446,  
18'd3958,  18'd12738,  18'd8997,  18'd2921,  -18'd13830,  -18'd3235,  
18'd17579,  18'd15364,  18'd12642,  -18'd2898,  -18'd5030,  18'd9907,  
18'd2023,  -18'd3024,  18'd6736,  18'd1395,  18'd4051,  18'd10703,  
-18'd33749,  -18'd11437,  -18'd25215,  18'd13106,  -18'd5154,  -18'd1430,  
-18'd21755,  -18'd1993,  -18'd2338,  18'd54162,  18'd13292,  18'd69454,  
18'd14556,  18'd19301,  18'd21515,  -18'd40546,  -18'd4808,  -18'd9132,  
-18'd16363,  18'd32247,  18'd15064,  18'd20156,  18'd10754,  18'd34371,  
-18'd5471,  -18'd4763,  18'd5134,  18'd3567,  -18'd2105,  18'd4521,  
18'd8828,  18'd19061,  18'd24016,  18'd16137,  -18'd15449,  18'd19753,  
18'd9486,  -18'd29362,  -18'd13787,  -18'd34336,  18'd11319,  -18'd8709,  
18'd2724,  18'd10420,  18'd12127,  18'd7352,  -18'd1843,  18'd33372,  


18'd15584,  18'd6919,  18'd1558,  -18'd14535,  -18'd3366,  -18'd9656,  
18'd13943,  18'd19863,  18'd23001,  -18'd58,  -18'd6547,  -18'd17828,  
-18'd17629,  18'd1657,  -18'd30530,  18'd19332,  18'd11198,  18'd15365,  
-18'd6625,  -18'd17627,  -18'd4547,  18'd9055,  -18'd5559,  18'd4957,  
-18'd1009,  18'd3010,  -18'd1716,  -18'd3352,  18'd443,  18'd3211,  
-18'd14484,  -18'd2020,  -18'd7751,  18'd15377,  18'd63,  18'd22578,  
-18'd5426,  18'd1800,  18'd12137,  -18'd24623,  -18'd316,  18'd7059,  
-18'd8017,  -18'd3068,  18'd8188,  18'd13251,  -18'd1885,  -18'd16474,  
-18'd18826,  -18'd1797,  -18'd14795,  18'd3960,  18'd6831,  18'd2384,  
-18'd11961,  -18'd15715,  -18'd4400,  18'd10394,  -18'd4412,  -18'd20307,  
-18'd4685,  -18'd37441,  18'd3367,  18'd5033,  -18'd7337,  18'd3495,  
-18'd7230,  18'd2570,  18'd6660,  18'd9309,  18'd175,  -18'd8575,  
-18'd1023,  18'd332,  -18'd3071,  -18'd7021,  18'd5613,  18'd1357,  
-18'd5478,  18'd12821,  18'd20073,  18'd29409,  -18'd5043,  18'd21947,  
-18'd9145,  -18'd8285,  -18'd10576,  -18'd10129,  18'd7787,  -18'd8902,  
18'd9697,  18'd10655,  -18'd3068,  18'd11903,  18'd8217,  18'd50,  

18'd2486,  18'd15422,  18'd12471,  18'd11541,  -18'd1519,  18'd3298,  
18'd11159,  18'd19890,  18'd22154,  18'd11587,  -18'd4054,  -18'd7108,  
18'd14513,  18'd14902,  -18'd27454,  -18'd17238,  18'd7240,  -18'd25919,  
18'd3079,  18'd8415,  18'd9724,  18'd20368,  18'd2361,  18'd33091,  
-18'd255,  -18'd82,  -18'd7733,  -18'd6161,  -18'd5558,  -18'd2439,  
-18'd11308,  -18'd20828,  -18'd27368,  18'd25350,  18'd4181,  18'd21064,  
-18'd26070,  -18'd39224,  -18'd17076,  18'd2242,  18'd11924,  18'd9919,  
-18'd1491,  18'd7052,  18'd13814,  18'd10064,  -18'd8879,  -18'd33052,  
18'd8928,  -18'd6446,  -18'd23491,  18'd10179,  18'd7603,  -18'd31899,  
-18'd13345,  -18'd27846,  -18'd1515,  -18'd21348,  18'd7338,  -18'd33083,  
-18'd3388,  -18'd10084,  18'd9809,  18'd14285,  18'd7298,  18'd12918,  
-18'd10817,  18'd15555,  -18'd4082,  18'd6266,  -18'd2309,  18'd876,  
-18'd6811,  -18'd7541,  18'd2337,  18'd3617,  -18'd440,  -18'd8497,  
18'd8001,  -18'd2925,  18'd797,  18'd19227,  -18'd8803,  18'd29982,  
-18'd3917,  -18'd14021,  -18'd16940,  -18'd25550,  18'd11130,  -18'd26010,  
18'd6805,  18'd7819,  18'd3834,  -18'd20364,  -18'd4423,  -18'd5837,  

-18'd18775,  -18'd28830,  -18'd19838,  18'd11564,  18'd3867,  -18'd7359,  
-18'd6312,  18'd122,  18'd22055,  18'd7207,  -18'd5359,  18'd8989,  
18'd21312,  18'd15484,  18'd12000,  -18'd56679,  -18'd3837,  -18'd36060,  
-18'd9230,  -18'd4117,  18'd9840,  18'd12275,  -18'd1082,  18'd9923,  
18'd1090,  18'd2522,  -18'd8622,  18'd4601,  18'd6111,  -18'd5271,  
18'd21681,  -18'd5096,  18'd3855,  -18'd2357,  -18'd2152,  -18'd21644,  
-18'd5743,  -18'd19299,  -18'd38065,  18'd5994,  18'd9419,  -18'd950,  
-18'd15024,  -18'd13965,  18'd18124,  -18'd3131,  -18'd5044,  -18'd17609,  
18'd22541,  18'd22030,  18'd19036,  -18'd17496,  -18'd14361,  -18'd3915,  
18'd9106,  -18'd3842,  18'd12073,  -18'd20522,  18'd3548,  18'd8851,  
18'd7625,  18'd7621,  -18'd6727,  -18'd8670,  18'd2706,  -18'd28691,  
18'd6292,  -18'd5923,  -18'd258,  18'd12522,  -18'd8423,  -18'd19244,  
-18'd629,  18'd3778,  -18'd4366,  -18'd1406,  -18'd94,  -18'd5983,  
-18'd2303,  18'd28446,  18'd16896,  18'd13257,  -18'd404,  18'd24701,  
-18'd4465,  -18'd8879,  -18'd2032,  -18'd25956,  18'd3076,  -18'd12358,  
18'd7470,  18'd10617,  -18'd8888,  -18'd4128,  18'd1815,  18'd13002,  

18'd2284,  -18'd7232,  -18'd6682,  -18'd22787,  -18'd2758,  -18'd29407,  
18'd5394,  -18'd5744,  18'd7405,  18'd20843,  -18'd11770,  18'd16815,  
18'd19231,  18'd29991,  18'd20565,  18'd3683,  -18'd13305,  18'd512,  
-18'd18681,  -18'd16864,  18'd12551,  18'd23274,  -18'd1863,  18'd18676,  
18'd5743,  -18'd6025,  18'd530,  18'd4072,  -18'd1848,  18'd3253,  
18'd14536,  18'd16826,  18'd22536,  18'd1323,  -18'd8423,  -18'd16800,  
18'd25167,  18'd13164,  -18'd10928,  -18'd29914,  18'd10379,  -18'd21951,  
-18'd3726,  -18'd24692,  18'd11557,  18'd14718,  18'd5339,  18'd2249,  
-18'd23356,  18'd3231,  18'd19623,  18'd32393,  -18'd1103,  18'd14634,  
-18'd10470,  18'd14714,  18'd2925,  18'd44098,  18'd3400,  18'd48336,  
18'd24796,  18'd12856,  18'd7927,  -18'd19509,  18'd2965,  -18'd45943,  
18'd15731,  18'd9126,  18'd18166,  -18'd4085,  -18'd9464,  -18'd16225,  
-18'd1504,  -18'd7309,  -18'd7536,  18'd539,  18'd5228,  -18'd7016,  
18'd4191,  18'd1602,  18'd555,  18'd14766,  -18'd10414,  18'd9477,  
-18'd1709,  -18'd18225,  -18'd13955,  -18'd16271,  18'd13160,  -18'd16571,  
-18'd15193,  -18'd19109,  -18'd33876,  -18'd9418,  -18'd1842,  18'd12238,  

18'd6470,  18'd19340,  18'd2799,  -18'd4693,  18'd1844,  -18'd8634,  
-18'd10919,  -18'd5825,  18'd20869,  18'd14638,  -18'd11613,  18'd10652,  
18'd891,  18'd4474,  18'd17447,  18'd13747,  -18'd6847,  -18'd6348,  
-18'd6325,  -18'd22871,  18'd9611,  18'd29471,  18'd5429,  18'd20876,  
-18'd4625,  -18'd1005,  18'd3632,  -18'd4034,  -18'd4642,  18'd5348,  
18'd12623,  18'd7267,  18'd29426,  18'd3970,  -18'd14658,  -18'd5290,  
18'd14944,  18'd26268,  18'd15101,  -18'd17959,  18'd7248,  18'd5984,  
-18'd3581,  18'd1803,  18'd15000,  18'd19860,  18'd2561,  18'd21580,  
-18'd32236,  -18'd37493,  -18'd30247,  18'd2516,  18'd4461,  -18'd22933,  
-18'd21847,  -18'd19728,  -18'd20265,  18'd40535,  18'd16984,  18'd34966,  
18'd1515,  18'd23542,  18'd18630,  -18'd15823,  -18'd5232,  18'd11678,  
-18'd45387,  -18'd4992,  18'd10250,  18'd30786,  18'd8687,  18'd25183,  
-18'd1034,  -18'd3885,  18'd1216,  18'd1737,  -18'd5093,  18'd4459,  
18'd9355,  18'd29539,  18'd28147,  -18'd543,  -18'd12590,  18'd11371,  
18'd5127,  -18'd19271,  -18'd5153,  -18'd42373,  18'd10454,  -18'd36643,  
-18'd10399,  18'd828,  -18'd29307,  -18'd2264,  18'd5777,  18'd27181,  


18'd18027,  18'd8287,  -18'd5388,  -18'd16695,  -18'd8036,  -18'd13760,  
18'd11389,  18'd20945,  18'd27296,  18'd22000,  -18'd6817,  18'd7933,  
-18'd2961,  -18'd1877,  -18'd9555,  18'd18217,  18'd9968,  -18'd10855,  
-18'd25327,  -18'd20982,  -18'd12027,  18'd27817,  18'd6361,  18'd11017,  
-18'd6236,  -18'd182,  18'd3353,  -18'd975,  18'd4212,  -18'd161,  
-18'd19335,  -18'd7942,  -18'd3963,  18'd8723,  -18'd5645,  18'd14436,  
-18'd8060,  -18'd1356,  18'd25468,  18'd108,  -18'd3984,  18'd18915,  
18'd2410,  18'd681,  18'd33672,  18'd24014,  -18'd9537,  18'd4369,  
-18'd9557,  -18'd2604,  18'd6358,  18'd23151,  -18'd5103,  18'd6989,  
-18'd13313,  -18'd18875,  -18'd16972,  -18'd18066,  -18'd7178,  -18'd14717,  
-18'd6077,  -18'd16212,  18'd424,  18'd6946,  18'd772,  -18'd161,  
-18'd4940,  18'd1967,  -18'd8205,  -18'd7756,  -18'd4552,  -18'd2309,  
-18'd4788,  18'd1507,  -18'd3648,  -18'd7432,  -18'd1097,  -18'd5772,  
-18'd3662,  18'd20443,  18'd29032,  18'd33316,  -18'd8349,  18'd31242,  
-18'd2730,  -18'd17414,  -18'd13435,  -18'd3958,  18'd7281,  -18'd15138,  
18'd16438,  18'd17054,  -18'd810,  18'd3411,  18'd2230,  18'd4563,  

-18'd41,  18'd18726,  18'd21416,  18'd8915,  -18'd2503,  -18'd3934,  
-18'd9957,  18'd3147,  18'd14330,  18'd24351,  -18'd4098,  18'd17478,  
18'd25936,  18'd13067,  18'd28138,  -18'd15285,  -18'd6866,  -18'd63042,  
18'd350,  18'd9717,  -18'd16142,  -18'd10285,  -18'd278,  18'd2969,  
18'd4852,  -18'd7168,  18'd3812,  18'd2782,  18'd2802,  18'd6482,  
-18'd13082,  -18'd10588,  18'd4411,  -18'd6106,  18'd5253,  18'd4367,  
-18'd32034,  -18'd32682,  -18'd35149,  18'd31683,  18'd9973,  18'd22659,  
-18'd966,  18'd5266,  18'd20636,  18'd16634,  -18'd7227,  18'd16918,  
-18'd56,  -18'd6697,  -18'd16170,  -18'd1126,  -18'd6613,  -18'd40485,  
-18'd7802,  -18'd26301,  18'd22142,  -18'd13127,  -18'd7833,  -18'd22780,  
-18'd20261,  -18'd8147,  -18'd11545,  18'd19085,  18'd5212,  18'd7334,  
-18'd1129,  18'd3913,  18'd1540,  18'd5547,  -18'd10359,  18'd1097,  
-18'd1894,  18'd580,  -18'd3054,  -18'd1584,  18'd5141,  -18'd6536,  
-18'd7617,  -18'd10833,  -18'd39516,  18'd29750,  -18'd6133,  18'd10985,  
-18'd4291,  -18'd7898,  18'd2446,  -18'd4405,  18'd4115,  -18'd22793,  
18'd11719,  18'd9536,  18'd11901,  -18'd3273,  -18'd1300,  18'd6585,  

-18'd10680,  -18'd29355,  -18'd4583,  18'd12186,  18'd3457,  -18'd12397,  
-18'd17500,  18'd449,  18'd2390,  18'd21695,  -18'd6399,  18'd24902,  
18'd22370,  18'd19912,  18'd36152,  -18'd2390,  -18'd2053,  18'd4897,  
18'd9932,  18'd11845,  18'd4275,  18'd1835,  -18'd3639,  18'd9796,  
-18'd1666,  -18'd4855,  -18'd4451,  18'd2173,  -18'd2111,  18'd1854,  
18'd12397,  -18'd8437,  -18'd13903,  -18'd20477,  -18'd6014,  -18'd16809,  
18'd8295,  -18'd13282,  -18'd34362,  18'd2180,  18'd14997,  -18'd5068,  
-18'd18058,  -18'd15600,  18'd8607,  18'd28983,  18'd2500,  18'd18753,  
18'd29693,  18'd24461,  18'd12871,  -18'd27312,  -18'd1745,  18'd4699,  
-18'd26408,  -18'd22897,  -18'd6301,  18'd28951,  18'd3455,  18'd6597,  
18'd14311,  18'd6111,  18'd2438,  18'd6548,  18'd4442,  -18'd22617,  
-18'd8684,  -18'd23846,  18'd21501,  -18'd7834,  -18'd4679,  -18'd11384,  
-18'd4523,  -18'd138,  18'd3396,  -18'd283,  -18'd4653,  -18'd2161,  
-18'd2883,  18'd34912,  -18'd5643,  18'd1003,  -18'd1536,  18'd18928,  
18'd2865,  -18'd8666,  -18'd5763,  -18'd6217,  18'd14147,  -18'd9208,  
18'd2168,  18'd3758,  18'd5174,  18'd10112,  18'd552,  18'd18640,  

-18'd1494,  -18'd15356,  18'd6083,  18'd5056,  18'd830,  -18'd24783,  
-18'd18039,  -18'd20200,  -18'd15591,  18'd15149,  18'd2943,  18'd19130,  
18'd6382,  18'd18214,  18'd16186,  18'd18449,  18'd839,  18'd6614,  
-18'd4694,  18'd13694,  18'd8177,  18'd8758,  18'd6320,  18'd11644,  
18'd1845,  -18'd1560,  -18'd6641,  -18'd1487,  -18'd5904,  18'd2882,  
18'd25547,  18'd15078,  18'd15856,  -18'd16469,  -18'd16950,  -18'd2237,  
18'd30802,  18'd25157,  18'd6092,  -18'd57797,  18'd9392,  -18'd35993,  
-18'd24645,  -18'd23149,  18'd4359,  18'd20238,  -18'd3723,  18'd26123,  
-18'd21507,  -18'd3718,  -18'd7054,  18'd17738,  18'd539,  18'd25040,  
-18'd7522,  -18'd3035,  -18'd14540,  18'd10872,  18'd5811,  18'd20416,  
18'd16583,  18'd19801,  18'd23467,  -18'd6307,  -18'd9458,  -18'd24506,  
-18'd6775,  18'd2251,  18'd2727,  18'd12623,  18'd1917,  18'd19956,  
18'd4080,  -18'd8076,  -18'd5930,  -18'd6816,  -18'd5708,  18'd5729,  
18'd5139,  -18'd2463,  -18'd14218,  18'd5452,  -18'd869,  18'd25305,  
18'd2118,  -18'd3570,  -18'd15444,  -18'd5419,  18'd4668,  -18'd15824,  
-18'd11249,  -18'd14763,  -18'd8865,  -18'd3497,  18'd6862,  18'd4990,  

18'd12610,  18'd5556,  -18'd3803,  -18'd16509,  -18'd6568,  -18'd7826,  
-18'd12918,  18'd613,  -18'd708,  18'd4710,  -18'd1485,  18'd19161,  
18'd20767,  18'd17802,  18'd13991,  18'd6688,  -18'd2110,  -18'd1450,  
-18'd6911,  18'd9101,  18'd2396,  18'd18250,  -18'd6522,  18'd4178,  
-18'd1230,  -18'd4680,  -18'd1846,  18'd3308,  18'd3839,  -18'd6083,  
18'd13677,  18'd18769,  18'd21446,  18'd6927,  -18'd15513,  18'd6003,  
18'd12879,  18'd38009,  18'd27357,  -18'd2915,  18'd7333,  18'd880,  
-18'd16378,  -18'd4444,  18'd8064,  18'd6660,  18'd8757,  18'd13935,  
-18'd31578,  -18'd39515,  -18'd16748,  18'd6538,  18'd2874,  -18'd8418,  
18'd8474,  -18'd3270,  -18'd20183,  -18'd882,  18'd8858,  -18'd16658,  
-18'd25440,  18'd12761,  18'd7860,  18'd14541,  -18'd131,  18'd23026,  
-18'd27727,  -18'd16917,  -18'd16542,  18'd22493,  -18'd3329,  18'd22645,  
-18'd2170,  -18'd3135,  18'd2322,  -18'd1336,  -18'd6373,  18'd2038,  
18'd9175,  18'd18572,  18'd2855,  18'd1316,  -18'd877,  18'd9954,  
18'd15829,  18'd1908,  -18'd15372,  -18'd28137,  18'd6859,  -18'd28044,  
-18'd19129,  -18'd28972,  -18'd18643,  18'd4320,  18'd260,  18'd12806
	};
	
	always @(posedge clk) begin
		if (rstn == 0) begin
			qa <= 0;
		end
		else if (!cena) begin
			qa <= weight[aa];
		end
	end
	
endmodule



