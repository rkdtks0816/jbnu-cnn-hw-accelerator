`include "global.sv"
`include "timescale.sv"
module wieght_fc2_rom(
	input			clk,
	input			rstn,
	input	[11:0]	aa,
	input			cena,
	output reg		[`WDP_WEIGHT*`OUTPUT_NUM_FC1*`OUTPUT_NUM_FC2 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC2*`KERNEL_SIZEX_FC2*`KERNEL_SIZEY_FC2-1][0:`OUTPUT_NUM_FC2-1][0:`OUTPUT_NUM_FC1-1][`WDP_WEIGHT-1:0] weight	 = {
18'd7345,  -18'd9197,  18'd13725,  18'd11819,  18'd9626,  18'd15827,  18'd27188,  18'd21512,  18'd2526,  -18'd16567,  -18'd38638,  18'd11461,  -18'd11588,  -18'd4935,  18'd10997,  -18'd2269,  
18'd12056,  18'd11702,  18'd10399,  -18'd41418,  18'd10295,  -18'd337,  18'd13608,  -18'd14281,  18'd9197,  18'd985,  18'd8787,  -18'd15925,  -18'd2294,  -18'd32135,  18'd13906,  -18'd7010,  
-18'd19274,  18'd950,  18'd6403,  18'd4453,  18'd14716,  18'd11395,  18'd8776,  -18'd11303,  18'd23811,  18'd31033,  18'd12431,  18'd2702,  18'd9274,  18'd2182,  18'd13586,  -18'd8970,  
-18'd12574,  -18'd6067,  18'd5386,  -18'd20476,  -18'd5507,  -18'd17716,  -18'd7466,  18'd10393,  18'd18916,  -18'd11172,  18'd28270,  18'd8779,  18'd12439,  18'd6420,  18'd14167,  18'd14199,  

18'd8044,  18'd1577,  -18'd934,  18'd9081,  -18'd2620,  18'd6465,  18'd13192,  -18'd28569,  -18'd26454,  -18'd625,  18'd977,  -18'd12088,  -18'd21433,  18'd14272,  -18'd2180,  18'd11947,  
-18'd77,  -18'd7066,  18'd25010,  18'd24137,  -18'd791,  18'd2027,  -18'd11544,  -18'd2023,  -18'd364,  -18'd8245,  -18'd23682,  18'd6389,  -18'd5547,  18'd20560,  18'd13269,  18'd16730,  
18'd791,  18'd794,  -18'd9028,  -18'd3247,  18'd1837,  -18'd4521,  18'd6111,  18'd11757,  -18'd35737,  -18'd5950,  -18'd8900,  -18'd5765,  -18'd15273,  18'd15227,  -18'd10052,  18'd2632,  
18'd6543,  18'd15158,  -18'd9242,  18'd25722,  18'd16327,  -18'd8380,  18'd18004,  18'd8964,  18'd20675,  -18'd4888,  -18'd823,  -18'd12763,  -18'd6649,  18'd24681,  -18'd18993,  18'd23940,  

-18'd11100,  18'd5961,  18'd19647,  18'd17939,  18'd20742,  -18'd16206,  18'd30074,  18'd39716,  18'd3735,  -18'd21861,  -18'd320,  -18'd1251,  18'd5029,  18'd5799,  18'd36048,  18'd3349,  
-18'd15026,  -18'd6567,  -18'd19075,  18'd2940,  -18'd11464,  -18'd245,  -18'd13647,  18'd20038,  -18'd10276,  -18'd13006,  -18'd21391,  -18'd8732,  -18'd28264,  -18'd15061,  18'd15852,  -18'd98,  
-18'd13890,  -18'd12232,  -18'd2439,  18'd7673,  -18'd625,  18'd22339,  18'd15425,  -18'd20922,  -18'd4237,  -18'd19292,  -18'd12497,  18'd8475,  18'd10478,  18'd27433,  -18'd21406,  -18'd3389,  
18'd10903,  18'd15292,  18'd2910,  18'd12602,  -18'd2305,  -18'd6708,  18'd6346,  -18'd14933,  18'd22621,  18'd6719,  18'd601,  18'd11227,  18'd19993,  -18'd27854,  -18'd12571,  18'd5279,  

-18'd13079,  18'd14588,  18'd17499,  -18'd23798,  18'd16286,  -18'd4525,  18'd277,  18'd3720,  18'd13307,  18'd12614,  -18'd23812,  18'd6332,  -18'd18493,  18'd20695,  18'd16105,  18'd23067,  
-18'd6473,  18'd12488,  18'd8031,  -18'd14433,  18'd2774,  18'd6250,  18'd7990,  18'd21174,  18'd13217,  -18'd9096,  18'd13218,  18'd3720,  18'd35704,  -18'd4333,  -18'd601,  -18'd12344,  
18'd16994,  18'd10269,  -18'd26478,  18'd3300,  18'd4346,  18'd16197,  18'd13712,  -18'd16481,  18'd3946,  -18'd28098,  -18'd14778,  -18'd13387,  18'd6234,  -18'd7383,  -18'd18697,  -18'd10062,  
18'd21984,  -18'd9622,  18'd145,  18'd11628,  -18'd5887,  18'd14045,  -18'd14867,  18'd8404,  18'd16453,  -18'd3698,  18'd25633,  18'd14122,  18'd13789,  -18'd9384,  -18'd23757,  -18'd10316,  

18'd14850,  18'd9385,  18'd16974,  18'd14019,  18'd35570,  -18'd9490,  -18'd14114,  -18'd510,  18'd18065,  18'd729,  18'd40495,  18'd16280,  18'd30885,  -18'd24087,  18'd21833,  -18'd5651,  
18'd82,  -18'd25722,  -18'd20918,  -18'd13661,  18'd7491,  18'd11166,  -18'd12362,  18'd18009,  -18'd625,  18'd17436,  -18'd14429,  18'd30214,  -18'd10731,  18'd3208,  -18'd7068,  -18'd12447,  
-18'd7323,  -18'd3267,  18'd23946,  -18'd12523,  18'd6243,  -18'd10715,  -18'd16973,  18'd13182,  -18'd20503,  18'd21480,  18'd8302,  -18'd407,  18'd6343,  18'd4693,  18'd22526,  -18'd8570,  
-18'd3212,  -18'd8415,  18'd1893,  -18'd2872,  18'd23659,  -18'd10935,  -18'd10826,  18'd1223,  18'd30637,  18'd4591,  -18'd14247,  18'd3092,  -18'd8594,  18'd1467,  -18'd677,  18'd20171,  

-18'd8373,  18'd15009,  18'd23787,  18'd5207,  -18'd322,  -18'd11028,  -18'd9073,  -18'd1262,  18'd16359,  18'd11812,  -18'd47611,  18'd4315,  18'd26217,  -18'd8717,  18'd4638,  -18'd1809,  
18'd9177,  18'd10675,  -18'd13889,  -18'd14161,  18'd23089,  18'd312,  -18'd15623,  -18'd22990,  18'd15800,  -18'd17983,  -18'd17234,  18'd15394,  -18'd10051,  -18'd19227,  -18'd9147,  -18'd20085,  
18'd13734,  18'd9845,  18'd2160,  18'd2463,  -18'd17311,  -18'd23254,  18'd8189,  -18'd2113,  -18'd519,  18'd31813,  18'd11010,  18'd10755,  -18'd10549,  -18'd7730,  -18'd13343,  18'd11808,  
18'd14717,  18'd20590,  18'd13514,  18'd15856,  18'd10342,  18'd20886,  18'd7015,  18'd12507,  -18'd29001,  -18'd7053,  18'd424,  18'd33623,  18'd7140,  18'd21742,  18'd26012,  -18'd3937,  

-18'd2954,  -18'd7987,  -18'd5802,  18'd9593,  -18'd10645,  18'd11564,  18'd9321,  18'd15594,  18'd3916,  -18'd5801,  -18'd12058,  -18'd16029,  -18'd19873,  -18'd8053,  -18'd6574,  -18'd5888,  
18'd530,  -18'd10647,  -18'd8399,  18'd28634,  18'd12290,  -18'd1184,  -18'd3587,  -18'd8475,  18'd7836,  18'd1164,  18'd8058,  18'd1374,  -18'd12137,  18'd22937,  -18'd4307,  18'd9689,  
-18'd11792,  18'd8431,  18'd5079,  -18'd2672,  -18'd10566,  -18'd11188,  18'd15929,  18'd14290,  18'd5753,  18'd15192,  -18'd10775,  18'd11381,  18'd8617,  -18'd6198,  -18'd558,  -18'd10589,  
-18'd873,  18'd18900,  -18'd15911,  -18'd25396,  -18'd1987,  -18'd3155,  -18'd8941,  -18'd3932,  -18'd20872,  -18'd8330,  18'd11252,  -18'd9500,  18'd164,  18'd15204,  18'd15492,  -18'd17588,  

-18'd1700,  -18'd1436,  18'd3169,  -18'd15379,  -18'd8460,  18'd9691,  -18'd15397,  18'd3524,  18'd15194,  18'd24085,  18'd2104,  -18'd6716,  -18'd12680,  18'd22397,  18'd10588,  -18'd11860,  
-18'd7404,  18'd10507,  -18'd14573,  -18'd6821,  18'd27780,  -18'd1958,  -18'd4072,  -18'd28458,  18'd504,  -18'd5927,  18'd22910,  18'd1588,  -18'd4141,  -18'd4548,  -18'd7029,  18'd19739,  
-18'd11546,  18'd12759,  -18'd8668,  18'd6096,  18'd5647,  -18'd15205,  -18'd15257,  -18'd10017,  18'd28241,  -18'd13303,  18'd26117,  -18'd10100,  -18'd15819,  18'd19882,  -18'd12068,  -18'd5994,  
-18'd2067,  18'd2561,  -18'd2632,  18'd16609,  -18'd14844,  18'd15021,  18'd27550,  -18'd6690,  -18'd24489,  18'd3635,  18'd3529,  18'd21948,  -18'd5445,  18'd41141,  -18'd13754,  18'd10356,  

18'd9553,  18'd4671,  -18'd5554,  18'd7422,  18'd19119,  18'd910,  18'd11512,  -18'd2,  18'd3168,  18'd21121,  18'd22049,  18'd7696,  18'd17849,  -18'd7851,  18'd10078,  -18'd2125,  
18'd9207,  18'd19592,  18'd15639,  18'd3961,  18'd11979,  18'd10861,  -18'd15133,  18'd4121,  18'd1172,  18'd12588,  18'd14255,  18'd30125,  18'd12487,  -18'd4617,  -18'd990,  -18'd30249,  
-18'd4367,  -18'd926,  18'd938,  18'd6732,  -18'd20097,  18'd10897,  18'd8801,  18'd53,  18'd184,  -18'd18553,  18'd7756,  18'd1227,  18'd13540,  18'd3597,  -18'd2879,  18'd4545,  
-18'd3288,  -18'd35636,  -18'd4365,  18'd4482,  -18'd8718,  -18'd13361,  18'd4518,  18'd13808,  18'd12168,  18'd2032,  -18'd1744,  18'd21814,  -18'd19543,  -18'd9082,  18'd22537,  18'd6082,  

18'd8568,  18'd19465,  18'd23603,  -18'd29866,  -18'd6350,  18'd8996,  -18'd7788,  -18'd11736,  18'd24786,  18'd8430,  18'd455,  -18'd6414,  -18'd14989,  -18'd14994,  18'd15051,  18'd15185,  
-18'd1249,  -18'd20488,  18'd25980,  -18'd982,  18'd3253,  18'd5893,  18'd9197,  -18'd566,  -18'd6483,  -18'd11653,  18'd29698,  18'd18220,  18'd12569,  18'd6963,  18'd4852,  18'd1951,  
-18'd9607,  18'd10206,  -18'd23723,  -18'd9021,  -18'd2148,  -18'd16842,  -18'd15858,  18'd6994,  18'd19087,  18'd2159,  -18'd12957,  18'd394,  18'd8807,  18'd14842,  -18'd8864,  -18'd665,  
18'd13468,  18'd18205,  -18'd2428,  -18'd2792,  -18'd89,  18'd15607,  18'd10555,  -18'd10715,  18'd29448,  18'd3268,  18'd26210,  18'd18373,  18'd12172,  18'd21018,  -18'd17779,  18'd24179,  

-18'd1130,  -18'd16280,  -18'd3589,  -18'd10325,  18'd5625,  -18'd6089,  18'd10357,  -18'd14756,  -18'd14137,  -18'd18325,  18'd73,  18'd16152,  -18'd10696,  18'd24716,  -18'd25638,  -18'd27397,  
18'd11,  -18'd6193,  -18'd702,  18'd8344,  -18'd13980,  -18'd9510,  -18'd4014,  18'd8315,  -18'd15305,  18'd15985,  -18'd6990,  18'd13421,  18'd17550,  18'd6677,  18'd9221,  -18'd3893,  
-18'd9263,  -18'd2894,  18'd19051,  -18'd1544,  18'd343,  -18'd13635,  18'd15932,  -18'd3287,  -18'd7331,  -18'd6081,  -18'd5235,  -18'd2556,  18'd13148,  18'd22327,  -18'd1427,  -18'd3214,  
18'd24887,  18'd8098,  18'd7292,  18'd21532,  18'd13087,  18'd18649,  18'd25264,  -18'd13039,  18'd15711,  18'd2868,  -18'd13475,  18'd4215,  -18'd15965,  -18'd8851,  18'd24563,  -18'd13210,  

18'd14576,  -18'd6774,  -18'd6914,  -18'd2734,  18'd18471,  18'd9846,  18'd1660,  -18'd3339,  -18'd5510,  -18'd1843,  -18'd16947,  18'd13768,  18'd1438,  18'd14545,  -18'd8149,  18'd1822,  
18'd8757,  18'd34548,  18'd25956,  18'd29637,  -18'd14125,  -18'd1634,  18'd6382,  18'd5224,  -18'd10361,  -18'd2438,  18'd21213,  -18'd21017,  18'd916,  -18'd4184,  -18'd363,  -18'd16772,  
-18'd14812,  18'd10522,  18'd19308,  18'd14054,  18'd6143,  18'd1210,  18'd8922,  18'd8346,  18'd25244,  -18'd4669,  -18'd16520,  -18'd10087,  18'd133,  18'd10390,  -18'd16308,  18'd13206,  
-18'd11892,  -18'd5699,  -18'd8971,  -18'd19664,  18'd10251,  -18'd23568,  18'd15018,  18'd9369,  -18'd18084,  18'd11545,  -18'd10413,  -18'd14420,  18'd20909,  18'd31288,  18'd10713,  -18'd24958,  

18'd6559,  -18'd3488,  18'd9585,  18'd8482,  18'd25944,  -18'd2138,  -18'd21213,  18'd9031,  18'd11580,  -18'd13882,  -18'd3373,  -18'd9873,  18'd7765,  18'd24391,  -18'd21230,  -18'd8241,  
-18'd1148,  18'd24331,  18'd23143,  18'd1638,  -18'd12369,  18'd7938,  18'd6269,  -18'd18795,  -18'd1371,  -18'd11515,  18'd15211,  18'd1652,  18'd18327,  -18'd22777,  -18'd6944,  18'd14415,  
-18'd342,  -18'd11923,  18'd1412,  -18'd9772,  18'd9178,  -18'd14190,  -18'd17501,  18'd3546,  18'd913,  18'd31371,  18'd2657,  -18'd7236,  18'd1502,  -18'd10969,  18'd23645,  18'd21123,  
18'd19836,  -18'd19107,  18'd2408,  18'd20956,  18'd4669,  -18'd8922,  18'd12831,  18'd1352,  18'd20721,  -18'd12227,  -18'd27830,  18'd17081,  -18'd16157,  18'd26632,  18'd152,  18'd2710,  

18'd14259,  -18'd12553,  -18'd5155,  -18'd10570,  18'd12982,  -18'd3698,  18'd4559,  18'd4306,  18'd2764,  -18'd17738,  18'd11157,  -18'd15275,  18'd9415,  -18'd12356,  -18'd3795,  18'd11858,  
18'd11763,  -18'd17,  -18'd9745,  -18'd7491,  -18'd5890,  18'd7825,  18'd5643,  -18'd11131,  18'd8574,  -18'd6914,  -18'd10893,  -18'd9178,  -18'd4251,  -18'd11726,  18'd11077,  -18'd4532,  
18'd9602,  -18'd15605,  18'd12298,  -18'd11561,  18'd6162,  18'd12733,  -18'd13208,  18'd10942,  18'd1412,  -18'd3774,  -18'd9615,  18'd9699,  -18'd2975,  18'd4348,  -18'd5394,  -18'd10108,  
-18'd5768,  18'd2192,  -18'd6851,  18'd4768,  18'd8897,  18'd4702,  18'd7179,  18'd1012,  -18'd12623,  18'd8754,  -18'd10204,  -18'd5230,  18'd383,  -18'd8863,  18'd12436,  18'd10420,  

18'd3617,  18'd7376,  -18'd2798,  -18'd27611,  18'd17743,  18'd3048,  18'd23200,  -18'd24011,  18'd7307,  18'd8670,  18'd12234,  -18'd9960,  18'd13738,  18'd1721,  18'd6248,  18'd22708,  
-18'd7266,  -18'd18470,  -18'd34101,  18'd29656,  18'd23438,  -18'd5625,  18'd13113,  18'd848,  -18'd12977,  18'd12435,  -18'd11940,  -18'd16156,  -18'd24483,  18'd6364,  -18'd1418,  -18'd7369,  
18'd5309,  18'd10946,  18'd6828,  -18'd2654,  18'd15092,  18'd17826,  18'd28967,  18'd26776,  -18'd1639,  -18'd1702,  18'd27104,  18'd13592,  -18'd5480,  18'd18870,  -18'd4229,  18'd12382,  
18'd14608,  -18'd20288,  -18'd7668,  18'd15725,  18'd12539,  -18'd22198,  -18'd45,  18'd15975,  -18'd27828,  18'd1951,  18'd7194,  -18'd13040,  18'd15429,  18'd10847,  -18'd5804,  -18'd16813,  

-18'd15578,  -18'd22772,  18'd15573,  18'd36550,  -18'd24193,  18'd11554,  18'd23378,  18'd9358,  -18'd1950,  18'd8339,  18'd1889,  -18'd626,  18'd15784,  18'd20130,  -18'd12721,  -18'd34053,  
18'd12218,  18'd8440,  18'd12452,  18'd34033,  18'd18392,  18'd3532,  -18'd11396,  18'd29454,  18'd14874,  -18'd4576,  -18'd232,  -18'd25568,  -18'd10149,  -18'd21560,  -18'd13996,  -18'd5589,  
-18'd9150,  18'd9086,  -18'd12820,  18'd13308,  18'd8520,  18'd21812,  18'd6974,  -18'd20181,  -18'd2957,  -18'd24113,  18'd25395,  -18'd2831,  -18'd9054,  -18'd5893,  -18'd11616,  18'd3255,  
18'd10535,  -18'd41259,  -18'd9979,  18'd8128,  18'd1251,  -18'd10815,  18'd25360,  -18'd16834,  18'd3291,  -18'd9334,  18'd10956,  -18'd15418,  18'd20940,  18'd6283,  18'd14070,  -18'd8086,  

18'd10340,  -18'd6880,  -18'd15520,  18'd17247,  18'd21219,  18'd13201,  18'd20279,  18'd28509,  18'd2559,  -18'd14688,  -18'd19893,  -18'd11032,  18'd11521,  18'd17778,  -18'd7365,  -18'd4588,  
18'd6025,  18'd25175,  18'd16821,  -18'd14953,  -18'd1108,  18'd7021,  18'd11765,  -18'd8812,  18'd14189,  18'd4595,  -18'd24754,  -18'd1205,  -18'd6042,  -18'd17660,  -18'd8789,  18'd30282,  
18'd12341,  -18'd5979,  -18'd7288,  18'd25,  18'd16287,  18'd12573,  -18'd9883,  -18'd5087,  -18'd18662,  -18'd1290,  -18'd17577,  18'd12811,  18'd2869,  18'd4053,  18'd7230,  18'd9535,  
18'd15335,  18'd27285,  -18'd6950,  -18'd2129,  -18'd18001,  18'd21277,  -18'd13218,  18'd4077,  -18'd1570,  -18'd1386,  -18'd2678,  -18'd4751,  -18'd18751,  18'd735,  18'd2081,  -18'd5110,  

-18'd403,  18'd1690,  -18'd16761,  -18'd12166,  -18'd14884,  18'd13101,  18'd4262,  -18'd9453,  -18'd8978,  18'd1501,  -18'd17543,  -18'd1249,  18'd17322,  -18'd4800,  18'd5273,  -18'd4178,  
18'd11871,  -18'd9580,  -18'd1869,  -18'd5226,  18'd7934,  -18'd9424,  -18'd11387,  -18'd7494,  18'd12247,  18'd15359,  -18'd796,  -18'd4017,  -18'd5053,  18'd9240,  18'd11968,  -18'd22125,  
18'd6147,  -18'd6956,  -18'd3444,  -18'd15054,  -18'd705,  18'd12264,  -18'd3462,  -18'd11184,  -18'd3815,  18'd10744,  -18'd5423,  18'd9383,  18'd7546,  18'd4335,  -18'd8257,  -18'd1614,  
-18'd18079,  -18'd8120,  -18'd12788,  18'd12172,  18'd14727,  -18'd13362,  -18'd4483,  18'd864,  18'd215,  -18'd14127,  18'd2548,  -18'd8480,  -18'd15107,  -18'd16101,  18'd3690,  -18'd13342,  

18'd7260,  -18'd13303,  -18'd11814,  -18'd31419,  18'd12092,  -18'd2752,  -18'd11194,  18'd10960,  18'd15159,  -18'd17740,  -18'd29181,  18'd11279,  18'd2085,  18'd13024,  -18'd7261,  18'd12900,  
-18'd1148,  -18'd9304,  18'd19020,  -18'd40056,  -18'd13777,  -18'd12474,  18'd2462,  18'd23076,  -18'd1761,  -18'd6973,  18'd17537,  -18'd29831,  -18'd17053,  -18'd12553,  18'd1315,  18'd10955,  
18'd7542,  -18'd4618,  18'd16086,  18'd1224,  18'd5522,  18'd9618,  -18'd6176,  -18'd5384,  18'd574,  -18'd14877,  18'd8421,  18'd12415,  -18'd12120,  18'd5347,  -18'd6790,  18'd5863,  
18'd3549,  18'd6820,  18'd4436,  18'd25285,  18'd24617,  18'd11158,  -18'd15696,  18'd9442,  18'd15162,  18'd7564,  18'd22006,  18'd5400,  -18'd19112,  18'd3301,  -18'd14429,  18'd13392,  

-18'd2595,  -18'd14399,  -18'd12517,  18'd18324,  -18'd7900,  18'd7704,  -18'd853,  -18'd12171,  -18'd10484,  -18'd16273,  -18'd18562,  18'd5372,  18'd12002,  18'd2681,  18'd3770,  18'd14656,  
18'd9586,  18'd18789,  18'd16090,  -18'd11632,  18'd17885,  -18'd7581,  18'd1045,  -18'd12521,  -18'd12877,  -18'd4169,  18'd24355,  18'd9277,  -18'd18926,  -18'd3013,  -18'd4871,  18'd21462,  
-18'd3052,  18'd2788,  18'd9038,  -18'd13673,  18'd14903,  18'd9621,  -18'd7836,  -18'd13932,  18'd30323,  -18'd12159,  -18'd6813,  18'd10780,  18'd11892,  18'd21968,  18'd5685,  -18'd8249,  
-18'd9686,  18'd7676,  -18'd7444,  -18'd934,  18'd8023,  -18'd9805,  18'd15020,  -18'd1574,  -18'd9655,  18'd6168,  18'd9398,  -18'd19103,  18'd8905,  -18'd6050,  18'd12777,  18'd32574,  

18'd13086,  -18'd19699,  18'd16119,  -18'd7797,  -18'd16814,  18'd8940,  18'd7645,  -18'd16618,  18'd6888,  18'd13528,  -18'd10921,  -18'd13233,  -18'd20315,  18'd2097,  -18'd743,  18'd6090,  
18'd11669,  18'd3695,  -18'd18292,  18'd18104,  -18'd12265,  18'd4847,  18'd9204,  -18'd6824,  -18'd244,  -18'd5944,  -18'd3456,  -18'd6251,  18'd21147,  18'd4031,  -18'd1159,  18'd3100,  
18'd5354,  18'd13579,  18'd288,  18'd15862,  -18'd16270,  -18'd17519,  18'd3639,  18'd7842,  -18'd32670,  -18'd5225,  18'd2766,  18'd724,  18'd1468,  18'd1223,  18'd7401,  -18'd15410,  
-18'd4834,  -18'd1962,  -18'd15280,  18'd674,  -18'd4348,  18'd17100,  18'd13634,  18'd10910,  -18'd13756,  18'd5869,  -18'd916,  -18'd3183,  -18'd21561,  18'd14777,  -18'd26883,  18'd13489,  

-18'd4880,  18'd18128,  18'd1040,  -18'd344,  18'd3176,  -18'd1057,  18'd2126,  18'd34138,  18'd10214,  18'd1698,  18'd8908,  18'd15488,  -18'd13741,  18'd6875,  18'd11850,  18'd9025,  
18'd1493,  18'd3902,  18'd9932,  18'd28506,  18'd6648,  -18'd1672,  -18'd13522,  18'd6751,  18'd3685,  -18'd11714,  18'd15278,  -18'd22337,  -18'd2722,  -18'd186,  18'd6210,  18'd21133,  
-18'd12066,  18'd7167,  -18'd16984,  18'd4629,  -18'd13457,  -18'd8096,  -18'd27825,  -18'd20956,  18'd139,  18'd2574,  -18'd7769,  18'd15967,  -18'd2284,  -18'd7607,  -18'd12891,  -18'd1543,  
-18'd8396,  18'd24712,  18'd2817,  -18'd13560,  18'd9087,  -18'd17952,  18'd7985,  18'd1611,  18'd21811,  -18'd13015,  -18'd9151,  18'd10441,  18'd1322,  -18'd3639,  18'd10681,  -18'd11588,  

18'd5375,  -18'd8905,  -18'd4052,  -18'd9453,  -18'd17023,  18'd4482,  -18'd1077,  -18'd8182,  -18'd15933,  -18'd11198,  -18'd11777,  -18'd8124,  18'd0,  18'd18444,  18'd23018,  18'd5929,  
-18'd2734,  -18'd24821,  18'd13336,  18'd10432,  18'd7700,  -18'd15091,  18'd4812,  18'd16498,  18'd825,  -18'd11687,  -18'd11083,  -18'd4601,  -18'd6374,  18'd20773,  18'd15335,  18'd13717,  
18'd12718,  18'd8758,  18'd19636,  18'd14901,  -18'd14395,  18'd16767,  18'd9057,  18'd17473,  18'd1256,  18'd27287,  18'd7597,  -18'd12748,  -18'd12414,  18'd11664,  18'd4915,  -18'd5895,  
18'd9942,  -18'd757,  18'd18683,  18'd22964,  18'd19544,  18'd310,  -18'd10519,  18'd11047,  -18'd3473,  18'd14958,  -18'd16261,  -18'd11976,  -18'd14642,  -18'd6189,  18'd7973,  18'd1392,  

-18'd10797,  18'd17530,  -18'd15119,  -18'd12881,  -18'd12367,  18'd13187,  -18'd18176,  18'd10927,  18'd9554,  -18'd18439,  -18'd8454,  -18'd463,  18'd24648,  18'd20008,  -18'd1970,  18'd1343,  
-18'd10682,  18'd16440,  -18'd31163,  -18'd22537,  -18'd4648,  -18'd724,  -18'd11262,  -18'd21738,  18'd14418,  -18'd7454,  -18'd22695,  -18'd8994,  18'd2541,  18'd15099,  -18'd1788,  -18'd8757,  
-18'd930,  -18'd214,  18'd16903,  -18'd12985,  18'd11527,  -18'd289,  18'd8756,  -18'd5975,  18'd12842,  18'd27116,  -18'd4163,  18'd14785,  -18'd9372,  -18'd5265,  18'd11657,  -18'd9971,  
18'd6612,  18'd23454,  -18'd16766,  18'd1394,  18'd11883,  18'd15852,  18'd789,  18'd2507,  -18'd30006,  -18'd11539,  -18'd17378,  18'd45,  18'd12998,  -18'd25574,  18'd22011,  -18'd391,  

18'd10717,  -18'd9013,  18'd1501,  18'd22703,  18'd5856,  18'd11867,  -18'd3144,  -18'd3711,  18'd7248,  18'd14182,  -18'd20732,  -18'd2095,  18'd391,  -18'd14301,  18'd11447,  -18'd3498,  
-18'd6839,  18'd8343,  -18'd20834,  18'd17464,  18'd9966,  18'd4229,  18'd2821,  -18'd3708,  -18'd3114,  18'd7168,  -18'd34139,  -18'd26735,  18'd16830,  18'd4486,  18'd10449,  18'd13855,  
-18'd18150,  18'd12719,  18'd4293,  18'd6897,  18'd4039,  -18'd20756,  -18'd5438,  18'd27755,  18'd13335,  -18'd15188,  18'd10878,  18'd13390,  -18'd8417,  18'd10568,  18'd19257,  18'd7653,  
18'd12010,  -18'd22088,  -18'd10059,  -18'd7397,  18'd10477,  18'd18644,  18'd27451,  -18'd11939,  -18'd25783,  -18'd6156,  18'd22933,  -18'd31001,  -18'd11931,  18'd20338,  18'd23035,  -18'd1199,  

-18'd13897,  -18'd2619,  -18'd11849,  -18'd20638,  -18'd11345,  18'd9272,  18'd18735,  18'd931,  18'd5639,  -18'd7709,  18'd9886,  18'd3142,  -18'd8093,  18'd10246,  18'd6666,  18'd11527,  
18'd10092,  18'd16768,  18'd61507,  -18'd19282,  -18'd7760,  -18'd346,  18'd4821,  18'd2591,  -18'd2204,  18'd13924,  18'd8099,  18'd5509,  18'd35878,  18'd16068,  -18'd14729,  -18'd16638,  
-18'd14698,  18'd3973,  18'd9178,  -18'd7810,  -18'd3241,  -18'd4671,  18'd13583,  18'd11447,  -18'd16074,  -18'd3167,  18'd378,  18'd2748,  -18'd2153,  -18'd18697,  18'd24545,  18'd11603,  
18'd14668,  -18'd9353,  -18'd8791,  18'd11695,  -18'd12983,  -18'd703,  -18'd14585,  18'd13596,  18'd19174,  18'd7627,  18'd10173,  -18'd1026,  -18'd13246,  18'd22333,  18'd2298,  18'd3207,  

18'd11212,  -18'd26259,  18'd9721,  18'd15226,  18'd1590,  -18'd16128,  -18'd11233,  18'd21528,  -18'd4064,  18'd20672,  18'd11571,  -18'd15155,  -18'd6233,  -18'd5691,  18'd7195,  18'd11817,  
-18'd8780,  18'd34748,  -18'd25297,  18'd7847,  -18'd6742,  -18'd15769,  18'd3124,  18'd21259,  -18'd15432,  -18'd2542,  18'd33668,  -18'd8034,  -18'd1436,  18'd3520,  18'd2376,  -18'd28217,  
-18'd7703,  -18'd5876,  18'd7644,  18'd4942,  -18'd1536,  18'd72,  18'd20118,  18'd20314,  -18'd26688,  18'd14490,  18'd2363,  -18'd6256,  -18'd12683,  18'd15672,  -18'd570,  18'd12171,  
18'd8086,  18'd18792,  -18'd509,  18'd18580,  -18'd4804,  18'd11686,  -18'd18778,  18'd4911,  18'd17104,  18'd1832,  18'd15819,  18'd9363,  -18'd8674,  18'd8796,  18'd23505,  18'd17420,  

18'd2079,  -18'd2690,  -18'd589,  18'd24358,  18'd4698,  18'd10597,  -18'd16177,  18'd14883,  -18'd14620,  18'd12349,  18'd19326,  -18'd4687,  -18'd23093,  18'd14639,  18'd16989,  18'd2125,  
-18'd13812,  -18'd3602,  -18'd1397,  18'd29890,  18'd6055,  -18'd468,  -18'd8581,  18'd18376,  -18'd11209,  -18'd5026,  18'd29363,  -18'd2028,  18'd8484,  18'd18233,  18'd10158,  -18'd10348,  
-18'd8381,  -18'd6381,  -18'd29577,  -18'd6819,  18'd10318,  -18'd10436,  -18'd10987,  18'd17553,  18'd4200,  -18'd13780,  -18'd18213,  -18'd9025,  -18'd12445,  -18'd14781,  -18'd19290,  18'd11241,  
-18'd15331,  18'd25419,  -18'd1981,  18'd13663,  18'd16668,  18'd3621,  18'd3513,  -18'd3409,  18'd10289,  18'd13051,  18'd7811,  18'd15936,  18'd14605,  18'd16802,  18'd16870,  18'd13038,  

-18'd2786,  -18'd12585,  -18'd14736,  18'd24342,  -18'd9718,  18'd16131,  -18'd2054,  18'd1590,  -18'd7704,  18'd25431,  18'd29417,  -18'd13981,  18'd23340,  -18'd9312,  -18'd6040,  18'd4199,  
-18'd15279,  18'd2989,  -18'd7640,  18'd13746,  -18'd14818,  18'd6409,  18'd17489,  18'd9407,  18'd12552,  18'd11754,  18'd8424,  -18'd8004,  18'd3669,  18'd14849,  18'd2939,  18'd15879,  
-18'd11108,  -18'd6482,  -18'd2692,  18'd15103,  18'd8986,  18'd16554,  18'd10780,  18'd4746,  -18'd9273,  18'd9796,  18'd22991,  18'd7943,  18'd15031,  18'd2706,  -18'd11631,  18'd19025,  
18'd3333,  18'd15914,  -18'd6893,  18'd1389,  18'd15208,  18'd30055,  18'd6903,  -18'd11041,  -18'd119,  18'd11008,  -18'd13374,  18'd16965,  18'd19209,  18'd15001,  18'd4137,  18'd1722,  

18'd6415,  18'd3494,  -18'd15342,  18'd3913,  -18'd16315,  18'd1008,  -18'd13535,  18'd11309,  -18'd13462,  18'd2276,  18'd11647,  18'd4765,  -18'd11589,  -18'd150,  -18'd13803,  -18'd1638,  
18'd10979,  18'd12039,  18'd11694,  18'd6212,  -18'd1533,  -18'd4015,  18'd1169,  18'd4782,  -18'd2364,  -18'd13221,  -18'd13952,  18'd10815,  -18'd10384,  -18'd9137,  18'd14311,  18'd383,  
18'd1334,  18'd11220,  -18'd7179,  -18'd3556,  -18'd4966,  18'd10016,  18'd4898,  -18'd1738,  18'd9191,  -18'd3236,  -18'd13427,  -18'd12212,  18'd12872,  -18'd8207,  -18'd14275,  -18'd5732,  
-18'd10638,  -18'd5027,  18'd2689,  -18'd4426,  -18'd12155,  -18'd6414,  18'd14609,  18'd2310,  18'd2054,  18'd16374,  18'd1644,  -18'd275,  -18'd7720,  -18'd11720,  -18'd5236,  -18'd13609,  

-18'd3360,  -18'd8961,  -18'd5616,  18'd15697,  -18'd5694,  18'd14440,  -18'd28634,  -18'd1787,  -18'd22383,  18'd3062,  18'd2136,  -18'd7314,  18'd16404,  18'd19118,  18'd6672,  -18'd17478,  
18'd786,  -18'd14634,  18'd18033,  -18'd4312,  18'd7245,  18'd5839,  -18'd3794,  18'd11654,  -18'd1760,  -18'd3906,  -18'd8751,  18'd32538,  -18'd19062,  -18'd27907,  18'd14293,  -18'd31362,  
18'd15081,  18'd6557,  -18'd1448,  -18'd8465,  -18'd11734,  -18'd21842,  18'd13453,  18'd9702,  18'd1043,  -18'd750,  -18'd595,  18'd10960,  18'd3466,  -18'd19066,  -18'd18286,  -18'd2905,  
18'd17701,  18'd5009,  18'd9380,  18'd3376,  18'd15253,  18'd15282,  -18'd4041,  18'd12943,  -18'd516,  18'd1129,  18'd5707,  18'd8221,  -18'd8227,  -18'd40402,  -18'd10326,  -18'd138,  

18'd7360,  18'd13396,  18'd8595,  -18'd15418,  18'd25010,  -18'd15832,  18'd5306,  -18'd5783,  18'd17679,  -18'd5600,  18'd24952,  -18'd15279,  18'd18553,  18'd18523,  -18'd12616,  18'd679,  
-18'd4877,  -18'd1385,  -18'd15123,  18'd12321,  -18'd17081,  -18'd7534,  -18'd12794,  18'd18192,  -18'd2409,  18'd7427,  -18'd22947,  -18'd10876,  18'd4493,  18'd9881,  18'd6877,  18'd4700,  
18'd5309,  -18'd12426,  18'd23942,  -18'd5481,  18'd4455,  18'd4339,  -18'd8914,  -18'd24097,  18'd8773,  -18'd9256,  18'd9095,  -18'd1796,  -18'd15276,  -18'd11465,  -18'd17837,  18'd14029,  
18'd8802,  18'd21424,  -18'd7062,  -18'd17808,  18'd16510,  18'd90,  -18'd10052,  -18'd7191,  18'd13486,  18'd8303,  18'd5671,  -18'd1764,  18'd6118,  -18'd37367,  18'd18550,  -18'd21027
	};
	
	always @(posedge clk) begin
		if (rstn == 0) begin
			qa <= 0;
		end
		else if (!cena) begin
			qa <= weight[aa];
		end
	end
	
endmodule



