`include "global.sv"
`include "timescale.sv"
module wieght_fc1_rom(
	input			clk,
	input			rstn,
	input	[11:0]		aa,
	input			cena,
	output reg		[`WDP_WEIGHT*`OUTPUT_NUM_CONV2*`OUTPUT_NUM_FC1 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC1*`KERNEL_SIZE_FC1*`KERNEL_SIZE_FC1-1][0:`OUTPUT_NUM_FC1-1][0:`OUTPUT_NUM_CONV2-1][`WDP_WEIGHT-1:0] weight	 = {
18'd7241,  -18'd6543,  -18'd3374,  -18'd1723,  18'd8547,  18'd8180,  -18'd8954,  -18'd9335,  -18'd4056,  -18'd1709,  -18'd8757,  18'd643,  -18'd2392,  -18'd1567,  18'd5230,  -18'd4508,  
-18'd5573,  -18'd8490,  18'd3196,  -18'd9369,  -18'd8532,  18'd2075,  18'd5044,  -18'd674,  -18'd4609,  18'd888,  -18'd2969,  18'd2380,  18'd4701,  -18'd1587,  18'd3544,  -18'd956,  
18'd897,  -18'd9109,  18'd7487,  -18'd9384,  18'd1635,  -18'd5052,  -18'd6435,  -18'd9237,  -18'd7721,  -18'd7519,  18'd3964,  18'd3072,  -18'd761,  -18'd2694,  18'd2514,  -18'd896,  
18'd6918,  18'd6916,  -18'd4529,  18'd3689,  -18'd1641,  -18'd2328,  18'd7527,  -18'd5829,  -18'd9408,  18'd7585,  -18'd7180,  18'd3030,  -18'd8689,  -18'd4471,  18'd5905,  18'd7983,  
18'd3558,  -18'd5956,  -18'd5397,  18'd566,  18'd5624,  18'd6332,  18'd5709,  -18'd1402,  -18'd1963,  -18'd4147,  -18'd771,  18'd7229,  18'd8710,  18'd4588,  18'd6911,  -18'd6674,  
-18'd3109,  18'd1377,  -18'd4949,  -18'd4384,  -18'd3133,  18'd6865,  18'd6768,  -18'd6566,  -18'd8452,  -18'd3429,  -18'd6604,  -18'd6850,  -18'd4345,  -18'd8847,  -18'd9326,  -18'd8135,  
18'd4725,  18'd801,  18'd6392,  18'd7342,  -18'd2388,  -18'd8349,  -18'd1474,  18'd3737,  -18'd4129,  18'd1518,  18'd8223,  -18'd1640,  18'd4040,  18'd979,  18'd2952,  -18'd149,  
18'd2800,  -18'd2201,  18'd1613,  -18'd7776,  -18'd1277,  18'd490,  18'd4740,  -18'd2618,  18'd16,  18'd6143,  18'd4505,  -18'd9486,  18'd2540,  18'd6673,  18'd4341,  18'd3709,  
-18'd5205,  18'd6342,  18'd5593,  18'd225,  18'd1739,  -18'd7474,  -18'd5514,  -18'd9472,  18'd5383,  -18'd7378,  -18'd1263,  18'd2589,  -18'd6815,  -18'd1279,  18'd3854,  18'd7298,  
-18'd7681,  -18'd7719,  18'd5434,  18'd157,  -18'd4576,  -18'd7865,  -18'd2422,  -18'd8199,  -18'd8130,  -18'd8167,  -18'd4548,  18'd4053,  18'd6665,  18'd1873,  18'd565,  -18'd7248,  
18'd4359,  18'd6664,  -18'd5344,  -18'd2616,  18'd1962,  18'd753,  -18'd4381,  18'd4599,  18'd2356,  18'd5548,  18'd358,  -18'd2402,  -18'd6090,  -18'd8829,  -18'd4344,  -18'd3330,  
-18'd7241,  -18'd897,  -18'd6931,  -18'd5567,  -18'd1232,  -18'd2557,  -18'd6530,  18'd6553,  -18'd275,  18'd1203,  -18'd4815,  -18'd7098,  18'd1935,  18'd5340,  -18'd4755,  -18'd9312,  
18'd2873,  18'd7881,  -18'd336,  18'd837,  18'd2159,  18'd6350,  18'd4908,  -18'd2177,  -18'd1673,  -18'd7442,  -18'd9275,  -18'd5456,  18'd4075,  -18'd9051,  -18'd2856,  18'd4371,  
-18'd5639,  -18'd3653,  -18'd2796,  -18'd751,  18'd2237,  18'd7017,  -18'd5924,  18'd6156,  -18'd5930,  -18'd8099,  -18'd5874,  18'd7344,  18'd585,  18'd7154,  -18'd8960,  -18'd6067,  
18'd5702,  18'd452,  -18'd3719,  -18'd389,  -18'd4984,  -18'd9054,  -18'd3753,  -18'd5468,  -18'd2673,  18'd982,  18'd3743,  18'd2293,  -18'd847,  -18'd1136,  18'd7334,  -18'd6851,  
18'd75,  -18'd3997,  18'd1821,  -18'd19,  -18'd8158,  18'd8091,  -18'd4510,  18'd1819,  18'd5296,  -18'd8712,  -18'd9121,  -18'd6692,  18'd2355,  -18'd2968,  -18'd8878,  -18'd1733,  

18'd5090,  -18'd11779,  18'd206,  -18'd376,  18'd7267,  18'd14209,  -18'd3585,  -18'd5320,  18'd22921,  18'd35159,  18'd4168,  18'd20744,  -18'd1155,  18'd14487,  18'd3906,  -18'd1086,  
18'd15679,  -18'd4813,  -18'd9161,  18'd17002,  18'd2744,  -18'd77,  -18'd5582,  18'd2063,  -18'd7500,  -18'd6530,  18'd5530,  18'd5003,  18'd2871,  18'd13408,  18'd4323,  18'd7322,  
-18'd3169,  18'd8154,  -18'd13379,  18'd1387,  18'd8171,  18'd884,  -18'd15739,  18'd3359,  -18'd30607,  -18'd18119,  -18'd12555,  -18'd18168,  18'd1586,  18'd9258,  -18'd10613,  18'd3630,  
-18'd15844,  18'd2294,  -18'd6966,  -18'd1239,  -18'd3478,  -18'd6766,  -18'd13565,  18'd7289,  18'd637,  -18'd2015,  -18'd6492,  -18'd7246,  -18'd2284,  18'd11749,  -18'd4291,  18'd6279,  
18'd14854,  18'd1985,  18'd6789,  -18'd11216,  -18'd5738,  18'd3035,  -18'd1850,  -18'd2020,  18'd1411,  18'd3118,  18'd2005,  -18'd1957,  -18'd7985,  18'd183,  18'd4445,  18'd3548,  
18'd14923,  -18'd7754,  -18'd12759,  -18'd6299,  -18'd6112,  -18'd5069,  18'd4172,  18'd2822,  18'd5991,  -18'd6765,  18'd9990,  18'd5071,  18'd129,  -18'd4429,  18'd5313,  -18'd1357,  
18'd4913,  18'd7897,  -18'd868,  -18'd7994,  18'd1144,  18'd2735,  18'd21140,  18'd10152,  -18'd1910,  18'd8172,  -18'd6830,  -18'd8358,  18'd9086,  18'd10492,  18'd2917,  -18'd362,  
-18'd16227,  -18'd9431,  18'd7469,  18'd4557,  -18'd8439,  18'd8289,  -18'd8742,  -18'd20342,  -18'd3098,  18'd23369,  18'd7560,  -18'd10359,  -18'd6517,  18'd9101,  -18'd12889,  -18'd2123,  
18'd12755,  18'd1671,  -18'd2311,  18'd3381,  -18'd1349,  18'd3300,  18'd1522,  18'd4316,  18'd14588,  -18'd6973,  -18'd13338,  -18'd3538,  -18'd5593,  -18'd6820,  18'd8575,  18'd6965,  
18'd11842,  18'd4848,  -18'd4189,  18'd11112,  -18'd4750,  -18'd60,  18'd9152,  -18'd1939,  -18'd5929,  18'd9823,  -18'd1950,  -18'd4318,  -18'd2480,  18'd1622,  18'd10142,  -18'd928,  
18'd1180,  -18'd5971,  18'd20590,  18'd12956,  18'd6734,  18'd5427,  18'd12381,  18'd14849,  -18'd3897,  18'd342,  18'd12732,  -18'd4056,  -18'd960,  -18'd2425,  -18'd4316,  -18'd3461,  
-18'd13845,  18'd14915,  -18'd13,  -18'd22240,  -18'd8259,  18'd13006,  18'd6564,  -18'd2078,  18'd1011,  18'd15254,  18'd8351,  18'd20066,  18'd3821,  18'd4813,  -18'd3641,  18'd364,  
-18'd4755,  18'd59,  -18'd6342,  18'd19484,  -18'd8256,  -18'd7520,  18'd5565,  -18'd2822,  18'd3897,  -18'd989,  -18'd6236,  18'd489,  18'd4356,  -18'd6700,  18'd14413,  18'd14317,  
18'd12112,  -18'd9971,  -18'd12192,  18'd27980,  -18'd323,  -18'd11610,  18'd8013,  -18'd5729,  -18'd6584,  -18'd770,  -18'd7115,  -18'd3133,  -18'd3005,  -18'd13833,  18'd19127,  -18'd3403,  
-18'd4250,  18'd5958,  18'd22565,  -18'd264,  18'd529,  18'd4402,  18'd9542,  18'd20508,  -18'd4042,  -18'd6259,  18'd14628,  -18'd9195,  -18'd3918,  -18'd15247,  18'd17287,  -18'd8375,  
-18'd13438,  18'd19568,  18'd21637,  18'd1338,  -18'd7127,  18'd2388,  18'd11840,  18'd13610,  -18'd7708,  18'd2054,  18'd6608,  18'd2841,  -18'd2293,  18'd7506,  -18'd5790,  18'd9953,  

-18'd758,  18'd11249,  -18'd9246,  -18'd19334,  18'd3842,  18'd7024,  18'd12661,  18'd20833,  18'd25891,  18'd10315,  18'd2597,  -18'd4098,  18'd6990,  18'd5195,  -18'd4964,  18'd2138,  
18'd27776,  -18'd11383,  -18'd11470,  18'd35571,  -18'd6609,  18'd9708,  18'd458,  -18'd14532,  18'd6292,  18'd26199,  18'd15695,  18'd16818,  18'd1703,  18'd11023,  18'd1635,  18'd6512,  
18'd14060,  18'd7976,  18'd7847,  18'd2820,  18'd6560,  18'd246,  -18'd4909,  18'd12796,  18'd5336,  18'd4633,  18'd3251,  18'd17378,  18'd369,  18'd9568,  -18'd8404,  -18'd3671,  
-18'd11942,  18'd16751,  18'd13853,  18'd13452,  -18'd4396,  -18'd2070,  -18'd3602,  18'd15040,  18'd16400,  -18'd18710,  -18'd13095,  18'd11393,  18'd9754,  -18'd2940,  18'd4554,  -18'd17971,  
18'd16532,  -18'd973,  18'd8859,  -18'd12489,  -18'd6100,  18'd1573,  -18'd10889,  -18'd10386,  18'd3190,  -18'd15043,  -18'd12572,  -18'd11854,  18'd10747,  -18'd887,  18'd10242,  18'd5767,  
18'd15047,  -18'd12233,  -18'd3738,  -18'd12852,  -18'd2256,  18'd5031,  18'd1152,  -18'd16203,  18'd163,  18'd2624,  18'd9156,  18'd7090,  18'd2688,  18'd9559,  -18'd7244,  18'd2882,  
-18'd4971,  18'd8679,  -18'd9702,  18'd607,  -18'd7431,  18'd3908,  -18'd786,  -18'd8718,  -18'd4529,  -18'd10211,  18'd8746,  18'd12974,  -18'd5827,  18'd716,  18'd8907,  18'd14054,  
-18'd23960,  18'd22441,  -18'd10668,  18'd146,  18'd1205,  -18'd6754,  -18'd7607,  -18'd1591,  -18'd2053,  -18'd503,  -18'd4079,  -18'd4447,  -18'd2015,  18'd14574,  18'd1173,  -18'd4768,  
18'd5572,  -18'd3198,  -18'd3238,  -18'd2884,  -18'd3767,  18'd3373,  18'd1104,  -18'd13453,  18'd6886,  -18'd13089,  -18'd11131,  -18'd9511,  18'd5560,  -18'd10561,  18'd5204,  18'd20639,  
18'd16406,  -18'd7448,  -18'd7080,  -18'd6513,  18'd6065,  -18'd1662,  18'd13779,  18'd9476,  -18'd1513,  18'd10692,  -18'd4564,  -18'd9857,  18'd4782,  -18'd6875,  18'd127,  18'd11131,  
-18'd6080,  -18'd11439,  -18'd3904,  -18'd11030,  -18'd2344,  -18'd4679,  18'd3684,  -18'd6816,  18'd11109,  18'd3322,  18'd13601,  18'd13695,  -18'd1473,  -18'd1042,  18'd13009,  -18'd2188,  
18'd1098,  -18'd11091,  -18'd2698,  -18'd3865,  18'd6834,  -18'd2074,  18'd8310,  -18'd10043,  -18'd8086,  18'd7345,  18'd17715,  18'd13876,  -18'd2962,  -18'd2007,  -18'd1907,  18'd5061,  
-18'd9006,  -18'd596,  18'd5798,  18'd3674,  18'd7501,  -18'd4064,  -18'd6700,  -18'd382,  18'd8362,  -18'd12230,  -18'd5821,  -18'd8303,  18'd4817,  -18'd14181,  18'd42,  18'd6089,  
18'd7629,  -18'd10983,  18'd1933,  18'd9037,  -18'd1549,  18'd7277,  18'd514,  -18'd2696,  -18'd7440,  18'd143,  18'd4822,  18'd10916,  -18'd110,  -18'd3470,  -18'd4404,  -18'd975,  
-18'd12163,  -18'd81,  18'd7210,  -18'd3946,  -18'd2110,  -18'd8023,  -18'd14911,  18'd3101,  18'd9069,  18'd5073,  -18'd9092,  -18'd12609,  18'd3449,  -18'd7974,  -18'd371,  -18'd9390,  
18'd5278,  18'd2123,  -18'd2438,  18'd3488,  -18'd5207,  -18'd17324,  18'd8703,  18'd14719,  18'd862,  18'd1285,  18'd6413,  18'd8346,  -18'd2660,  -18'd6935,  18'd2967,  -18'd14583,  

-18'd39296,  -18'd10648,  -18'd16455,  18'd15320,  -18'd6926,  -18'd32384,  18'd3712,  18'd21008,  -18'd52818,  18'd1912,  -18'd3174,  -18'd14731,  18'd4256,  -18'd21936,  18'd2253,  -18'd20195,  
-18'd28583,  18'd8029,  18'd4608,  -18'd22651,  -18'd927,  -18'd2098,  18'd9083,  18'd16350,  -18'd48521,  -18'd904,  18'd6697,  -18'd6128,  -18'd5257,  18'd4214,  -18'd3334,  -18'd24348,  
-18'd22427,  18'd16163,  18'd17689,  -18'd5560,  18'd847,  18'd19249,  -18'd11059,  18'd11766,  18'd6197,  18'd31568,  18'd20497,  18'd7392,  18'd3132,  18'd733,  -18'd8976,  18'd5510,  
18'd16152,  -18'd4380,  -18'd17329,  18'd25323,  18'd1911,  -18'd379,  -18'd10323,  -18'd15016,  18'd14037,  18'd19257,  -18'd5898,  18'd12247,  18'd3199,  18'd11889,  18'd3677,  18'd27632,  
-18'd8375,  -18'd19192,  -18'd50,  18'd12423,  -18'd3445,  -18'd13023,  -18'd8568,  -18'd11929,  -18'd36512,  -18'd6427,  -18'd5297,  -18'd3396,  -18'd740,  -18'd11057,  18'd6638,  -18'd21704,  
-18'd5515,  -18'd3712,  18'd4735,  -18'd13982,  18'd5004,  18'd3666,  18'd12694,  -18'd1975,  -18'd9151,  -18'd2642,  18'd8239,  -18'd10488,  18'd4351,  -18'd3776,  18'd6679,  -18'd11689,  
-18'd16979,  18'd10021,  18'd15099,  -18'd12012,  18'd608,  18'd10522,  18'd9396,  18'd22928,  -18'd6387,  18'd2275,  -18'd14023,  -18'd14413,  18'd4541,  18'd12589,  18'd6314,  -18'd860,  
-18'd752,  -18'd3251,  -18'd7397,  18'd25346,  -18'd2576,  -18'd6044,  18'd7233,  -18'd5408,  18'd11352,  -18'd20901,  -18'd1697,  -18'd11800,  18'd8972,  18'd6339,  18'd4177,  -18'd1621,  
-18'd3593,  18'd9037,  -18'd11956,  18'd21021,  -18'd165,  -18'd13262,  -18'd2311,  18'd21604,  -18'd12005,  18'd7747,  18'd1517,  18'd1381,  18'd409,  -18'd6757,  -18'd2905,  -18'd14107,  
18'd4657,  -18'd8009,  18'd11080,  -18'd25468,  -18'd2486,  18'd6690,  18'd5696,  -18'd4633,  18'd2997,  18'd8852,  -18'd3524,  -18'd3510,  -18'd6202,  18'd2101,  18'd395,  -18'd7746,  
18'd2480,  18'd4847,  18'd9126,  -18'd10124,  -18'd6298,  18'd17694,  18'd3188,  18'd10293,  18'd10936,  -18'd8377,  -18'd11119,  -18'd8791,  -18'd3906,  18'd3374,  18'd2926,  18'd1121,  
18'd8783,  18'd22098,  -18'd6034,  18'd11493,  18'd4869,  18'd4616,  18'd14361,  18'd8697,  18'd207,  18'd6746,  -18'd3470,  -18'd4128,  -18'd1159,  -18'd1673,  -18'd4876,  18'd16028,  
-18'd11718,  18'd7177,  -18'd615,  18'd24895,  18'd5567,  18'd1898,  18'd6721,  -18'd10084,  -18'd21216,  -18'd2418,  18'd16487,  -18'd3556,  -18'd5712,  18'd7299,  -18'd5594,  -18'd9065,  
18'd12502,  -18'd5365,  -18'd1178,  -18'd5248,  -18'd1440,  18'd20717,  18'd9679,  -18'd1719,  18'd8612,  -18'd8504,  18'd14297,  -18'd129,  -18'd7813,  18'd9361,  -18'd3272,  -18'd8487,  
-18'd2488,  18'd5531,  18'd8058,  18'd16756,  18'd7070,  18'd6439,  -18'd6611,  18'd8226,  18'd13798,  -18'd4164,  -18'd6008,  -18'd7385,  18'd1692,  -18'd13775,  -18'd1810,  18'd15544,  
18'd18125,  18'd13007,  -18'd3670,  18'd19430,  -18'd5298,  -18'd13621,  18'd2151,  18'd18677,  -18'd5462,  18'd12208,  -18'd14827,  -18'd1148,  18'd4970,  -18'd2819,  18'd11421,  18'd9929,  

18'd10722,  18'd15645,  18'd9185,  18'd18727,  -18'd5561,  -18'd4528,  -18'd14849,  -18'd8141,  -18'd2907,  -18'd1757,  -18'd5592,  -18'd11643,  -18'd10375,  18'd12259,  -18'd7023,  18'd19563,  
18'd18560,  18'd571,  -18'd6847,  18'd9690,  18'd5886,  18'd1065,  -18'd14025,  18'd22343,  -18'd16919,  18'd6164,  18'd2078,  -18'd13211,  18'd3618,  18'd831,  18'd6721,  18'd1811,  
-18'd14247,  18'd724,  -18'd7645,  18'd20032,  -18'd6154,  -18'd7094,  -18'd13528,  18'd11668,  -18'd11502,  -18'd6405,  -18'd4395,  -18'd2728,  18'd4765,  -18'd4509,  18'd15181,  -18'd1614,  
-18'd9750,  18'd6750,  -18'd24489,  18'd2933,  18'd178,  -18'd14676,  -18'd12644,  18'd20603,  -18'd45744,  18'd1235,  18'd18204,  -18'd203,  18'd4370,  18'd5701,  18'd7667,  -18'd13024,  
18'd17096,  18'd8162,  -18'd3968,  -18'd3746,  18'd4740,  -18'd3289,  -18'd1039,  -18'd9712,  18'd4876,  18'd52,  -18'd10825,  -18'd11884,  -18'd10792,  -18'd967,  -18'd756,  18'd2374,  
18'd20123,  -18'd90,  -18'd915,  18'd4873,  -18'd4054,  -18'd3507,  18'd291,  -18'd2200,  -18'd388,  -18'd7684,  -18'd6534,  18'd7933,  -18'd8025,  -18'd3403,  18'd1199,  18'd4641,  
18'd8729,  18'd2257,  -18'd11614,  18'd5149,  -18'd5162,  18'd14039,  18'd14366,  18'd17507,  -18'd5572,  18'd9585,  -18'd4345,  -18'd1260,  18'd3116,  18'd4359,  18'd15523,  -18'd1974,  
-18'd5029,  18'd5096,  18'd24812,  -18'd4422,  -18'd8603,  18'd8409,  18'd15886,  -18'd14614,  -18'd24209,  18'd2150,  18'd27336,  -18'd1032,  -18'd3713,  18'd8767,  -18'd1221,  18'd4579,  
18'd26780,  18'd9471,  -18'd1920,  18'd8586,  18'd3347,  18'd16496,  18'd7608,  -18'd1785,  18'd1413,  -18'd25478,  -18'd10689,  -18'd2198,  -18'd7151,  -18'd4556,  -18'd1645,  18'd7408,  
18'd24034,  18'd8649,  -18'd4515,  18'd15067,  18'd6973,  -18'd9768,  -18'd1203,  -18'd3109,  18'd9039,  18'd8913,  18'd1064,  -18'd5147,  18'd1707,  18'd3965,  18'd7725,  18'd11727,  
18'd6012,  18'd4368,  18'd12905,  18'd10157,  -18'd6357,  -18'd3704,  -18'd2210,  18'd177,  18'd7013,  18'd9527,  18'd8584,  18'd8678,  -18'd6330,  -18'd9446,  18'd14459,  -18'd1184,  
18'd8672,  18'd15192,  18'd11686,  -18'd6137,  -18'd1764,  18'd19343,  18'd9658,  -18'd2002,  18'd5367,  18'd17587,  18'd10832,  18'd3624,  -18'd8457,  18'd16027,  18'd4304,  18'd11548,  
-18'd1121,  18'd5486,  18'd9425,  18'd15235,  -18'd605,  18'd6176,  18'd3129,  -18'd4296,  18'd8130,  -18'd23568,  -18'd8955,  -18'd25750,  -18'd3700,  18'd13562,  -18'd9573,  18'd24492,  
18'd8373,  18'd16719,  18'd2544,  18'd44436,  -18'd5872,  18'd3719,  18'd3941,  -18'd10673,  18'd3232,  -18'd542,  -18'd4504,  -18'd6799,  -18'd11220,  18'd3475,  -18'd1515,  18'd16723,  
-18'd2428,  18'd31683,  18'd3156,  18'd16463,  18'd3537,  -18'd16626,  -18'd9914,  18'd7548,  -18'd89,  18'd11484,  -18'd8267,  -18'd10035,  -18'd6958,  18'd64,  18'd2132,  18'd9697,  
-18'd10804,  18'd18800,  -18'd15715,  18'd439,  18'd1018,  -18'd5638,  18'd6372,  18'd23564,  -18'd9369,  18'd5251,  18'd8799,  -18'd6096,  -18'd3523,  18'd9343,  -18'd7089,  18'd4979,  

18'd3117,  18'd356,  18'd1063,  18'd6538,  18'd1523,  18'd278,  -18'd230,  -18'd11301,  -18'd1318,  -18'd7846,  -18'd6831,  -18'd4622,  -18'd2425,  18'd5258,  18'd6450,  -18'd5715,  
-18'd3385,  -18'd114,  18'd6382,  -18'd4785,  18'd6800,  -18'd2458,  -18'd5983,  -18'd4741,  -18'd3578,  18'd2199,  -18'd9560,  18'd172,  -18'd3739,  -18'd5937,  18'd2310,  -18'd5655,  
18'd5173,  -18'd3465,  -18'd1685,  18'd5351,  18'd4422,  -18'd5804,  18'd4037,  -18'd2759,  18'd3683,  -18'd10855,  -18'd2524,  -18'd11311,  18'd6840,  -18'd5973,  -18'd4903,  18'd3301,  
-18'd2237,  18'd7106,  -18'd6507,  -18'd7979,  18'd3748,  18'd524,  18'd668,  -18'd5628,  -18'd1274,  -18'd9551,  -18'd3372,  -18'd9601,  -18'd7821,  18'd373,  -18'd11115,  18'd1057,  
-18'd5384,  -18'd6877,  -18'd269,  18'd4133,  -18'd8062,  18'd2327,  -18'd1036,  18'd1680,  -18'd8918,  -18'd1655,  -18'd4508,  18'd6273,  18'd1986,  -18'd9342,  18'd2236,  18'd5852,  
-18'd1485,  -18'd11751,  -18'd7321,  18'd2703,  18'd1179,  -18'd6849,  -18'd6961,  18'd3330,  -18'd6746,  -18'd1102,  -18'd7202,  -18'd10157,  -18'd2174,  -18'd8547,  18'd460,  -18'd7177,  
-18'd1190,  18'd4346,  -18'd6711,  18'd1302,  18'd1640,  -18'd869,  18'd3180,  -18'd10970,  -18'd940,  -18'd2665,  -18'd5306,  18'd3984,  18'd8566,  -18'd6694,  18'd3347,  -18'd2803,  
18'd6300,  18'd6548,  18'd3179,  -18'd922,  -18'd2969,  18'd3121,  18'd3938,  18'd4986,  -18'd6711,  -18'd12327,  18'd4986,  -18'd9444,  18'd1179,  18'd2985,  18'd2819,  -18'd474,  
18'd1914,  -18'd300,  -18'd7699,  18'd2765,  -18'd3592,  18'd2863,  -18'd12009,  18'd4042,  -18'd5916,  -18'd6095,  18'd4677,  -18'd6075,  18'd3680,  18'd1448,  18'd1108,  18'd3581,  
18'd3981,  -18'd3131,  -18'd3171,  -18'd1617,  -18'd768,  -18'd415,  18'd1677,  -18'd9065,  -18'd2314,  18'd4676,  18'd1621,  18'd2274,  -18'd4803,  -18'd3068,  -18'd9588,  -18'd1790,  
18'd3970,  -18'd3100,  18'd5961,  18'd1921,  18'd1402,  -18'd1417,  18'd3033,  -18'd10348,  18'd4826,  -18'd8125,  18'd2494,  -18'd5905,  18'd2468,  -18'd4784,  -18'd1016,  18'd799,  
18'd6252,  -18'd1596,  18'd1019,  -18'd4502,  -18'd1254,  18'd478,  18'd760,  -18'd3026,  -18'd165,  -18'd4512,  18'd1769,  -18'd1291,  18'd4784,  -18'd6456,  18'd1150,  18'd7106,  
-18'd2601,  -18'd11148,  -18'd4519,  18'd2706,  18'd3744,  -18'd1985,  18'd4618,  -18'd1431,  -18'd1498,  -18'd5404,  18'd3982,  -18'd1004,  18'd200,  -18'd717,  -18'd201,  -18'd10353,  
18'd103,  18'd136,  -18'd2971,  18'd2739,  -18'd3999,  -18'd690,  -18'd4316,  18'd7168,  -18'd7368,  -18'd7192,  -18'd9768,  -18'd10447,  -18'd2245,  -18'd6532,  18'd4407,  18'd4604,  
-18'd4057,  18'd2267,  -18'd10330,  -18'd7369,  -18'd2935,  18'd1382,  -18'd5476,  -18'd5293,  18'd6016,  18'd3192,  -18'd131,  -18'd9484,  18'd2143,  18'd1318,  -18'd10721,  18'd7316,  
18'd4473,  -18'd4339,  18'd2985,  18'd5286,  -18'd5898,  -18'd8283,  -18'd6453,  -18'd6228,  -18'd7114,  18'd5039,  -18'd4479,  18'd487,  -18'd4236,  -18'd6250,  -18'd5381,  -18'd5470,  

18'd16329,  18'd1040,  18'd2181,  -18'd11763,  -18'd8018,  18'd4836,  -18'd9087,  -18'd488,  -18'd144,  18'd952,  -18'd15775,  18'd12260,  18'd5290,  18'd18843,  -18'd2897,  -18'd3469,  
18'd9047,  18'd176,  18'd1668,  18'd26377,  18'd4612,  -18'd8411,  18'd2739,  18'd335,  18'd4438,  18'd23835,  18'd7572,  -18'd2983,  18'd1392,  -18'd3990,  18'd10238,  -18'd10050,  
18'd9929,  -18'd15031,  18'd6911,  -18'd3668,  -18'd3740,  -18'd3849,  18'd7393,  18'd10236,  18'd12544,  18'd9706,  -18'd74,  18'd17705,  18'd8586,  -18'd13756,  18'd20462,  -18'd10012,  
-18'd4409,  -18'd6359,  18'd4304,  -18'd17262,  -18'd3990,  -18'd11362,  18'd10874,  18'd16988,  18'd22348,  -18'd12061,  18'd13134,  18'd21007,  18'd919,  -18'd6280,  18'd27786,  -18'd10588,  
18'd4725,  -18'd9431,  -18'd3234,  -18'd5368,  18'd8586,  -18'd8534,  18'd5208,  -18'd6062,  -18'd1244,  18'd7180,  18'd5146,  18'd4990,  18'd1058,  18'd3677,  18'd11973,  -18'd8772,  
18'd10656,  -18'd15595,  -18'd10007,  18'd7364,  18'd1480,  -18'd7423,  18'd1041,  -18'd20619,  -18'd4283,  18'd24772,  18'd6028,  18'd2708,  -18'd3985,  18'd4726,  18'd6982,  -18'd3818,  
-18'd3404,  -18'd4488,  -18'd11599,  18'd18301,  18'd3241,  -18'd11362,  -18'd11983,  18'd4757,  18'd3611,  18'd1667,  -18'd6121,  18'd7325,  -18'd5239,  18'd1870,  18'd11228,  -18'd12809,  
-18'd3206,  18'd652,  18'd10455,  -18'd5497,  -18'd8454,  -18'd3381,  18'd9736,  18'd13330,  -18'd15759,  -18'd32885,  18'd1644,  18'd5494,  18'd8265,  -18'd11536,  18'd18925,  18'd2788,  
-18'd1142,  18'd6204,  18'd11124,  -18'd11984,  18'd1787,  -18'd5703,  18'd9688,  -18'd1047,  -18'd1889,  -18'd362,  18'd1473,  18'd1564,  18'd8091,  18'd5621,  18'd3310,  -18'd800,  
18'd12149,  -18'd13081,  -18'd3043,  18'd6652,  18'd3118,  18'd9125,  18'd560,  -18'd250,  18'd5363,  18'd13079,  18'd2662,  18'd9463,  -18'd1093,  -18'd2162,  18'd5556,  18'd3122,  
18'd4843,  -18'd14129,  -18'd1928,  -18'd5433,  -18'd2079,  18'd10138,  -18'd18754,  18'd3831,  18'd1045,  18'd7040,  18'd1597,  18'd18013,  -18'd4624,  18'd10635,  18'd15474,  -18'd4526,  
18'd4041,  -18'd9254,  18'd13009,  -18'd2226,  18'd6003,  18'd2436,  18'd5436,  18'd12643,  -18'd1499,  -18'd20182,  -18'd7817,  18'd3163,  18'd1104,  18'd5511,  -18'd1130,  -18'd2875,  
18'd13612,  18'd4730,  18'd9683,  -18'd3937,  18'd6810,  18'd7044,  18'd1928,  18'd18484,  18'd2549,  -18'd2801,  18'd2806,  -18'd8905,  -18'd6091,  18'd2147,  -18'd1724,  18'd2645,  
18'd10655,  18'd1895,  18'd7891,  18'd7957,  -18'd5156,  18'd1947,  -18'd1825,  18'd13574,  -18'd5527,  18'd10462,  -18'd5746,  -18'd1066,  18'd2027,  18'd5830,  -18'd5232,  -18'd11418,  
-18'd5916,  18'd16205,  18'd4504,  18'd11213,  18'd4593,  18'd4355,  -18'd23325,  18'd5108,  -18'd7112,  18'd2675,  18'd4835,  18'd18193,  18'd11525,  18'd8132,  -18'd7865,  18'd6611,  
18'd3575,  18'd7035,  -18'd12764,  -18'd4269,  18'd866,  -18'd9724,  -18'd16007,  18'd9597,  -18'd7488,  -18'd7200,  18'd6081,  18'd7162,  18'd6734,  18'd7398,  -18'd3993,  -18'd13259,  

-18'd5053,  -18'd1075,  18'd7698,  -18'd4519,  -18'd8367,  18'd8743,  -18'd4836,  -18'd6213,  18'd22964,  -18'd10507,  18'd5860,  -18'd788,  -18'd8981,  18'd2240,  18'd966,  18'd26894,  
-18'd4454,  18'd5671,  18'd2247,  18'd9292,  -18'd8822,  18'd1789,  -18'd3830,  18'd8538,  -18'd6375,  -18'd1982,  -18'd481,  -18'd12009,  18'd399,  18'd4387,  -18'd6602,  18'd23059,  
-18'd7431,  18'd16127,  -18'd5500,  18'd2827,  -18'd6829,  -18'd1727,  18'd17164,  18'd6185,  -18'd553,  -18'd4837,  18'd7472,  -18'd10343,  18'd2114,  18'd648,  -18'd3652,  18'd11380,  
-18'd224,  18'd10452,  18'd10872,  18'd9241,  18'd7622,  18'd3387,  18'd16079,  18'd6279,  -18'd26719,  18'd9254,  -18'd2982,  18'd10977,  18'd234,  -18'd5948,  -18'd18031,  -18'd9219,  
18'd3424,  18'd18758,  18'd343,  -18'd3694,  18'd3053,  18'd16562,  18'd5041,  -18'd3289,  18'd6148,  -18'd10381,  18'd5367,  18'd10287,  -18'd6814,  18'd14060,  -18'd13062,  18'd10825,  
18'd5444,  18'd1965,  18'd4323,  18'd9145,  18'd109,  -18'd6793,  -18'd23225,  -18'd10704,  18'd8064,  -18'd274,  -18'd2443,  -18'd7961,  18'd2167,  -18'd6972,  -18'd12185,  18'd11621,  
18'd15489,  -18'd6560,  18'd5825,  -18'd6849,  -18'd7038,  -18'd9214,  18'd426,  18'd11192,  -18'd3589,  -18'd877,  18'd6692,  -18'd7122,  -18'd6574,  -18'd11938,  18'd5912,  18'd7867,  
-18'd623,  -18'd8301,  18'd17000,  -18'd2949,  18'd2578,  18'd17726,  -18'd43,  18'd4111,  18'd11730,  18'd21263,  18'd13157,  18'd10700,  -18'd2331,  -18'd4351,  18'd5422,  -18'd15565,  
18'd18652,  18'd10437,  18'd17833,  18'd21094,  18'd2779,  18'd5623,  18'd1507,  -18'd13106,  -18'd619,  -18'd21454,  18'd11443,  18'd3885,  18'd1732,  18'd12728,  -18'd9286,  18'd11018,  
-18'd9240,  -18'd2183,  -18'd7691,  -18'd6299,  -18'd7442,  18'd164,  -18'd18487,  -18'd6114,  -18'd2361,  18'd4725,  -18'd24277,  -18'd17694,  -18'd11103,  18'd1034,  -18'd11050,  18'd202,  
18'd10760,  -18'd4057,  -18'd23819,  18'd9204,  -18'd9145,  -18'd13815,  -18'd4169,  18'd17469,  -18'd6086,  -18'd2044,  18'd435,  -18'd5366,  18'd1512,  -18'd16367,  -18'd6514,  -18'd2318,  
18'd315,  18'd6522,  -18'd15538,  -18'd5239,  -18'd2375,  18'd1763,  18'd12128,  18'd17645,  18'd4611,  18'd8636,  18'd13860,  18'd3925,  18'd1146,  18'd4338,  -18'd6684,  -18'd8418,  
-18'd1940,  -18'd439,  18'd13140,  -18'd12051,  -18'd4015,  18'd7535,  -18'd10924,  -18'd17992,  18'd8859,  -18'd34076,  -18'd10667,  -18'd9448,  -18'd2877,  18'd12909,  -18'd9394,  18'd19722,  
-18'd8408,  -18'd6134,  18'd9639,  -18'd4142,  -18'd1081,  -18'd4922,  -18'd30353,  -18'd5295,  18'd2860,  18'd11906,  -18'd13806,  -18'd6022,  -18'd9658,  -18'd6792,  -18'd13588,  18'd15658,  
-18'd5084,  -18'd11254,  -18'd25081,  18'd17790,  18'd305,  -18'd33731,  -18'd17315,  -18'd6653,  -18'd20872,  18'd13666,  -18'd13759,  -18'd11099,  18'd6328,  -18'd16210,  18'd4791,  -18'd11365,  
-18'd19593,  -18'd12097,  -18'd25155,  18'd220,  -18'd2527,  -18'd14547,  18'd14665,  18'd7319,  -18'd15532,  18'd4882,  -18'd204,  18'd6636,  -18'd557,  -18'd11272,  18'd438,  -18'd38532,  

18'd27329,  -18'd15537,  18'd4952,  -18'd20880,  18'd1609,  18'd20158,  18'd5952,  -18'd8106,  18'd29863,  18'd13189,  18'd5343,  18'd27458,  -18'd5059,  18'd7219,  18'd12502,  18'd2086,  
18'd25291,  -18'd16182,  -18'd5695,  18'd2683,  18'd4954,  18'd8613,  -18'd12185,  18'd1820,  18'd18720,  18'd4470,  18'd4616,  18'd774,  18'd6920,  18'd7926,  -18'd304,  18'd7370,  
18'd3169,  18'd2835,  -18'd10757,  18'd726,  -18'd6712,  -18'd23625,  -18'd13674,  18'd9230,  -18'd22369,  18'd5961,  -18'd11909,  -18'd13212,  -18'd6801,  -18'd2436,  -18'd12386,  -18'd2796,  
-18'd28958,  18'd8775,  -18'd10593,  18'd12505,  -18'd3799,  -18'd9186,  -18'd18576,  18'd18638,  -18'd18380,  18'd10294,  -18'd1623,  -18'd991,  18'd2157,  18'd107,  -18'd20256,  -18'd7215,  
18'd31495,  18'd8099,  18'd5105,  -18'd31997,  18'd5951,  18'd11365,  -18'd2384,  18'd3336,  18'd8102,  -18'd13032,  -18'd3175,  18'd4176,  18'd8713,  18'd2413,  18'd781,  18'd8332,  
18'd6485,  18'd2845,  18'd143,  -18'd24622,  -18'd3774,  18'd1260,  18'd8588,  18'd4526,  18'd17899,  -18'd1796,  18'd9570,  18'd5612,  18'd7072,  -18'd5399,  -18'd6440,  -18'd4074,  
18'd15656,  -18'd10499,  18'd1718,  -18'd2384,  18'd8317,  -18'd8063,  18'd7906,  18'd5484,  18'd7220,  18'd18420,  18'd9228,  18'd11317,  18'd2155,  -18'd9123,  18'd1874,  -18'd325,  
-18'd2374,  18'd7323,  -18'd13783,  18'd2790,  -18'd6206,  18'd13083,  -18'd4223,  -18'd17286,  -18'd2366,  18'd31830,  -18'd1858,  18'd6063,  18'd408,  18'd16715,  -18'd1625,  -18'd3158,  
18'd230,  -18'd6713,  18'd4686,  -18'd15717,  -18'd1490,  18'd3795,  18'd8990,  18'd1806,  18'd13611,  -18'd12633,  -18'd1813,  -18'd243,  -18'd3981,  -18'd17797,  -18'd4131,  18'd22506,  
-18'd1572,  18'd7942,  -18'd10141,  18'd3163,  18'd408,  18'd3966,  18'd18645,  18'd1687,  18'd6022,  18'd7768,  -18'd7920,  -18'd10293,  -18'd7683,  -18'd2505,  18'd11526,  18'd13608,  
-18'd1568,  -18'd12014,  18'd11016,  18'd5765,  18'd3377,  -18'd6556,  18'd12696,  -18'd13522,  -18'd911,  18'd12957,  -18'd1060,  18'd5124,  -18'd879,  -18'd18933,  18'd4668,  -18'd3531,  
18'd6682,  -18'd10752,  -18'd3780,  -18'd14576,  -18'd5899,  18'd2806,  18'd13568,  -18'd14202,  18'd2188,  18'd3051,  18'd15252,  18'd17084,  18'd8734,  18'd6451,  18'd6779,  -18'd12700,  
-18'd16263,  18'd4140,  18'd8524,  -18'd432,  -18'd2973,  18'd3583,  18'd3188,  18'd3395,  18'd14854,  18'd6917,  -18'd14429,  -18'd1344,  18'd6485,  -18'd2222,  -18'd2484,  18'd23257,  
18'd13018,  18'd3563,  -18'd7878,  18'd11594,  -18'd6815,  -18'd5884,  -18'd7977,  -18'd4593,  18'd8045,  18'd7613,  -18'd9527,  -18'd5234,  18'd4971,  -18'd2282,  18'd11984,  18'd16548,  
-18'd9289,  -18'd6828,  18'd8277,  18'd2506,  -18'd1844,  18'd1955,  18'd4223,  18'd14365,  18'd3383,  18'd6794,  18'd11202,  -18'd13160,  18'd6628,  -18'd14598,  -18'd5268,  -18'd1236,  
-18'd17403,  18'd21,  18'd1925,  -18'd3147,  18'd2851,  -18'd14710,  18'd16158,  18'd13788,  -18'd20656,  18'd7723,  18'd10965,  18'd2306,  18'd5758,  -18'd13261,  18'd6852,  -18'd5076,  

-18'd2456,  -18'd14138,  18'd19260,  -18'd5463,  -18'd8047,  18'd2095,  18'd1795,  18'd7089,  18'd11829,  18'd442,  -18'd3187,  18'd8160,  18'd5078,  -18'd6110,  18'd11494,  -18'd21171,  
-18'd10846,  -18'd15271,  -18'd1907,  18'd7112,  18'd5231,  18'd5109,  -18'd7679,  -18'd4757,  18'd10037,  18'd4642,  -18'd8985,  18'd26909,  18'd9469,  18'd21388,  18'd1039,  -18'd19554,  
18'd1742,  18'd3211,  -18'd5521,  18'd14667,  18'd1169,  18'd10655,  -18'd8078,  -18'd5308,  -18'd2371,  18'd6338,  -18'd7056,  18'd8811,  18'd6521,  18'd14284,  -18'd11846,  18'd3914,  
18'd2143,  18'd10917,  -18'd8546,  -18'd246,  18'd8348,  18'd21957,  -18'd3239,  18'd19049,  18'd8576,  -18'd8808,  -18'd21656,  18'd12423,  18'd10221,  18'd8391,  -18'd2867,  18'd5686,  
18'd2131,  18'd13967,  18'd4294,  18'd1396,  18'd5133,  -18'd1941,  -18'd8618,  18'd11073,  -18'd11914,  -18'd19534,  18'd6324,  -18'd389,  -18'd5520,  -18'd6279,  18'd4857,  18'd7936,  
18'd556,  18'd5822,  -18'd4396,  -18'd8563,  -18'd1922,  -18'd11885,  18'd7856,  18'd4308,  -18'd9616,  -18'd8821,  -18'd14311,  -18'd11622,  18'd6177,  18'd14388,  18'd11890,  -18'd8735,  
-18'd3380,  -18'd11643,  18'd644,  18'd5840,  18'd4420,  18'd1355,  -18'd5532,  -18'd2878,  -18'd3764,  18'd4803,  -18'd7996,  -18'd12850,  18'd3530,  18'd3674,  -18'd153,  -18'd14720,  
18'd16582,  18'd4646,  18'd2538,  18'd7322,  -18'd3411,  18'd981,  -18'd9536,  18'd6277,  18'd18766,  18'd5862,  18'd8969,  18'd11485,  18'd3222,  18'd3816,  18'd2074,  -18'd11875,  
-18'd8969,  -18'd3316,  -18'd5286,  -18'd4909,  -18'd8076,  18'd6328,  18'd625,  18'd4384,  -18'd1380,  -18'd2308,  -18'd3041,  -18'd2965,  18'd1116,  -18'd5469,  -18'd4600,  18'd7769,  
-18'd11027,  -18'd11483,  18'd6312,  -18'd27678,  -18'd1209,  -18'd3468,  -18'd6578,  -18'd6428,  -18'd9402,  18'd2602,  18'd318,  -18'd384,  18'd4830,  -18'd4398,  18'd5327,  18'd4347,  
18'd9274,  18'd5706,  -18'd7400,  -18'd10178,  18'd5884,  18'd3528,  18'd13848,  18'd414,  -18'd3807,  -18'd811,  -18'd1360,  -18'd7576,  18'd10677,  18'd7752,  18'd1023,  -18'd7255,  
18'd7632,  18'd9696,  18'd9778,  18'd524,  18'd4873,  18'd10759,  -18'd2878,  18'd660,  18'd453,  18'd5067,  18'd10023,  -18'd3859,  18'd3102,  18'd3975,  18'd9026,  -18'd805,  
18'd6275,  18'd1246,  18'd6296,  -18'd11545,  -18'd2022,  18'd8046,  18'd12489,  18'd1107,  -18'd13848,  -18'd2261,  -18'd5802,  -18'd2605,  18'd8917,  -18'd4865,  18'd349,  18'd5561,  
18'd1809,  -18'd16127,  18'd14256,  -18'd29791,  -18'd5580,  18'd5381,  18'd2505,  18'd4371,  -18'd2430,  18'd5304,  18'd15124,  -18'd1082,  -18'd4605,  -18'd12905,  18'd11762,  18'd10067,  
18'd9180,  -18'd11552,  18'd1784,  -18'd14292,  18'd6440,  18'd6576,  -18'd1351,  18'd6663,  18'd16308,  18'd4804,  -18'd1481,  18'd1674,  18'd408,  18'd1267,  18'd12486,  18'd8525,  
-18'd1629,  18'd18294,  18'd9030,  -18'd7147,  -18'd2709,  18'd2787,  18'd13959,  18'd1348,  18'd8920,  18'd4837,  18'd4361,  -18'd7756,  18'd5351,  -18'd3298,  -18'd3849,  -18'd1442,  

-18'd5868,  18'd20623,  18'd10733,  -18'd5751,  -18'd5221,  18'd6991,  -18'd4791,  18'd12998,  18'd1902,  18'd2783,  18'd9165,  18'd19387,  -18'd6015,  18'd4481,  18'd1860,  -18'd5629,  
-18'd11432,  18'd2579,  -18'd2087,  -18'd14705,  -18'd7903,  -18'd11553,  -18'd854,  18'd1385,  -18'd4392,  -18'd16499,  -18'd8506,  -18'd9780,  -18'd7375,  18'd13253,  -18'd4552,  18'd3747,  
-18'd18236,  18'd1432,  -18'd10529,  18'd23463,  18'd1574,  18'd2650,  -18'd17320,  -18'd9227,  -18'd1143,  -18'd6284,  -18'd7269,  -18'd1736,  -18'd9357,  -18'd11625,  -18'd14728,  -18'd14952,  
18'd17563,  18'd3959,  -18'd32730,  18'd507,  18'd464,  18'd4793,  18'd986,  18'd6868,  18'd7727,  -18'd18541,  -18'd16018,  18'd117,  18'd5056,  18'd3804,  -18'd15255,  -18'd29546,  
18'd3914,  -18'd2430,  18'd2538,  -18'd7889,  -18'd6226,  18'd5708,  -18'd2220,  18'd2127,  -18'd1669,  -18'd1601,  -18'd1979,  18'd4786,  18'd2694,  18'd5624,  -18'd8416,  18'd3159,  
18'd11486,  18'd4741,  18'd121,  18'd888,  -18'd2951,  -18'd15553,  -18'd9179,  18'd3454,  18'd2666,  -18'd2359,  18'd2139,  -18'd10468,  -18'd3696,  18'd9989,  18'd3538,  18'd1898,  
-18'd9789,  18'd15996,  18'd10756,  -18'd5583,  -18'd4721,  -18'd136,  -18'd22561,  18'd5312,  18'd4291,  18'd2952,  18'd17073,  -18'd12399,  -18'd381,  18'd8737,  -18'd7714,  -18'd748,  
18'd2676,  18'd5698,  -18'd4185,  18'd2078,  -18'd4834,  -18'd2804,  -18'd18202,  -18'd6522,  -18'd4789,  18'd13645,  -18'd21606,  -18'd4608,  -18'd58,  -18'd1770,  -18'd26987,  18'd10892,  
-18'd11326,  18'd801,  18'd3131,  -18'd9802,  -18'd6224,  18'd13112,  -18'd1689,  18'd1380,  18'd8208,  -18'd14789,  18'd5876,  18'd9727,  -18'd7198,  18'd966,  18'd2561,  -18'd9010,  
18'd8573,  -18'd5193,  -18'd482,  -18'd13840,  -18'd6465,  18'd501,  -18'd10478,  -18'd19078,  18'd3570,  -18'd8839,  18'd9790,  18'd7923,  -18'd6528,  18'd1087,  -18'd1506,  18'd3078,  
18'd421,  18'd21383,  18'd8786,  -18'd6275,  -18'd126,  18'd12594,  18'd8389,  18'd9544,  18'd8042,  18'd2474,  18'd8778,  18'd3026,  -18'd8050,  -18'd4934,  18'd5521,  18'd10684,  
18'd10841,  18'd5691,  18'd9579,  18'd16303,  -18'd7118,  -18'd20250,  18'd5756,  -18'd25719,  18'd4530,  18'd18315,  -18'd1296,  18'd432,  18'd3331,  18'd1381,  18'd14685,  18'd19172,  
18'd3020,  18'd1349,  18'd8598,  -18'd32712,  18'd29,  18'd7195,  18'd12121,  18'd1357,  18'd13986,  -18'd19008,  18'd2489,  18'd9204,  18'd2240,  18'd1886,  -18'd13605,  18'd1491,  
-18'd9941,  18'd9873,  18'd15112,  -18'd7424,  -18'd2319,  18'd8630,  -18'd5064,  18'd3561,  18'd4073,  18'd1163,  -18'd7605,  -18'd2390,  -18'd7594,  -18'd2499,  -18'd9978,  18'd11194,  
18'd6532,  18'd5741,  18'd13830,  18'd11717,  -18'd5766,  -18'd18383,  -18'd14842,  -18'd6553,  18'd13019,  -18'd2774,  -18'd7257,  -18'd9298,  -18'd6534,  18'd404,  18'd2803,  18'd11214,  
-18'd13961,  18'd4905,  -18'd10426,  -18'd1360,  18'd8136,  -18'd28296,  18'd6594,  -18'd13580,  -18'd20547,  -18'd7202,  18'd9634,  -18'd11964,  -18'd1610,  -18'd8690,  18'd10794,  18'd9560,  

-18'd6494,  18'd5342,  -18'd7337,  -18'd900,  18'd1512,  -18'd10077,  -18'd4080,  18'd3795,  -18'd3388,  -18'd6186,  -18'd1788,  18'd1698,  18'd7997,  18'd4014,  18'd3703,  18'd3915,  
18'd2698,  18'd2706,  -18'd6822,  -18'd1415,  -18'd2553,  18'd200,  -18'd9121,  18'd1628,  -18'd6061,  18'd717,  18'd2842,  18'd2819,  18'd6644,  18'd5511,  -18'd8275,  -18'd9718,  
-18'd1709,  18'd8142,  -18'd6890,  18'd4990,  18'd6086,  -18'd4096,  18'd1949,  18'd60,  18'd855,  -18'd119,  -18'd9953,  -18'd7563,  18'd385,  18'd3201,  18'd6006,  18'd2246,  
-18'd1680,  -18'd3291,  -18'd8596,  -18'd1760,  -18'd7972,  18'd1668,  -18'd3953,  18'd8396,  -18'd2855,  18'd6918,  -18'd4612,  -18'd5555,  18'd5189,  -18'd8231,  18'd4466,  -18'd408,  
-18'd500,  18'd4107,  -18'd359,  18'd6657,  -18'd4006,  -18'd818,  18'd5544,  -18'd9061,  18'd3792,  -18'd8657,  18'd5352,  18'd6138,  18'd3463,  18'd458,  18'd2278,  18'd8104,  
-18'd2161,  18'd8368,  18'd2977,  -18'd8580,  -18'd5515,  -18'd820,  18'd4506,  -18'd8038,  -18'd3737,  -18'd920,  -18'd1891,  18'd3778,  18'd5535,  18'd5610,  -18'd320,  -18'd5275,  
-18'd3152,  18'd2013,  18'd5353,  -18'd8842,  -18'd4273,  -18'd6667,  -18'd3697,  -18'd3674,  18'd2219,  -18'd1845,  -18'd6637,  18'd576,  -18'd1215,  18'd4536,  -18'd6843,  -18'd5823,  
18'd5508,  -18'd7718,  -18'd2344,  18'd5898,  18'd5611,  18'd1048,  -18'd1736,  -18'd8149,  18'd1816,  -18'd5392,  18'd4584,  18'd650,  18'd920,  18'd4107,  -18'd3796,  -18'd3257,  
-18'd7495,  -18'd2995,  -18'd7175,  18'd3313,  18'd7523,  -18'd3728,  18'd3846,  18'd823,  18'd1401,  18'd4953,  -18'd8331,  18'd2275,  -18'd675,  -18'd3681,  -18'd2443,  -18'd6576,  
18'd4560,  -18'd7026,  -18'd5421,  -18'd450,  -18'd4316,  -18'd8791,  -18'd4062,  18'd2277,  -18'd5486,  18'd2572,  -18'd3920,  18'd5074,  -18'd523,  -18'd8760,  18'd1293,  18'd1559,  
-18'd7823,  -18'd9626,  -18'd1911,  -18'd1634,  -18'd2435,  -18'd2629,  18'd663,  18'd3663,  18'd1498,  18'd3798,  18'd2774,  -18'd4684,  -18'd4705,  18'd2341,  -18'd6695,  18'd3911,  
-18'd9501,  18'd4489,  -18'd769,  -18'd9520,  -18'd4054,  -18'd810,  -18'd8825,  -18'd4761,  -18'd7752,  -18'd490,  -18'd7677,  -18'd5989,  18'd4494,  -18'd6326,  -18'd9325,  18'd3506,  
18'd6185,  -18'd2892,  18'd6381,  -18'd7444,  18'd6609,  -18'd6359,  -18'd196,  18'd2958,  -18'd7459,  18'd5677,  -18'd3408,  18'd5908,  -18'd4470,  -18'd7602,  18'd6666,  -18'd944,  
-18'd10583,  18'd2493,  -18'd2493,  -18'd2825,  18'd7262,  -18'd2261,  18'd4486,  18'd4164,  -18'd10105,  -18'd6271,  -18'd7607,  18'd2006,  18'd7320,  -18'd6653,  -18'd5769,  18'd3941,  
-18'd6122,  18'd3939,  18'd5817,  18'd3492,  -18'd4457,  -18'd4951,  -18'd7336,  -18'd2713,  -18'd9517,  18'd2498,  18'd8683,  18'd5267,  18'd1962,  -18'd7231,  18'd1371,  -18'd5072,  
-18'd10107,  -18'd1868,  18'd1291,  -18'd9592,  -18'd6419,  18'd4559,  -18'd2854,  -18'd5439,  -18'd5224,  18'd4822,  -18'd8911,  -18'd9728,  18'd2730,  18'd5709,  -18'd5738,  -18'd8596,  

-18'd8405,  -18'd2469,  -18'd11978,  -18'd4745,  -18'd7063,  -18'd5525,  -18'd6203,  18'd6867,  -18'd10562,  18'd17778,  18'd6287,  18'd23085,  18'd5009,  -18'd82,  18'd14636,  -18'd21984,  
-18'd1026,  -18'd11433,  18'd3335,  -18'd17437,  18'd4686,  18'd11877,  -18'd9805,  18'd1921,  18'd5495,  18'd13789,  -18'd6996,  18'd9537,  18'd2568,  18'd12077,  -18'd1769,  -18'd4089,  
18'd3331,  -18'd12029,  18'd293,  -18'd429,  -18'd6470,  18'd6060,  -18'd16602,  18'd8708,  -18'd3631,  18'd14499,  18'd21009,  -18'd4893,  -18'd4006,  18'd1149,  18'd5470,  18'd5830,  
18'd14018,  18'd996,  -18'd6005,  18'd18139,  18'd6426,  -18'd12954,  -18'd28777,  18'd4500,  -18'd6499,  18'd24455,  18'd20541,  18'd11397,  -18'd6133,  18'd427,  18'd3897,  18'd17625,  
18'd10114,  18'd8785,  -18'd11263,  -18'd28798,  18'd5631,  -18'd7433,  18'd3481,  18'd15674,  -18'd20490,  18'd3356,  18'd11101,  -18'd5523,  18'd5947,  -18'd4571,  18'd13424,  -18'd1582,  
-18'd3173,  -18'd4860,  18'd5934,  -18'd10759,  -18'd6424,  18'd2809,  18'd12421,  18'd4743,  18'd6758,  -18'd13936,  18'd8553,  -18'd7596,  -18'd1561,  18'd390,  18'd5905,  -18'd9020,  
18'd1596,  18'd5106,  18'd16200,  -18'd5949,  18'd6623,  18'd17355,  18'd30207,  18'd3490,  18'd6852,  -18'd6632,  -18'd3293,  -18'd13096,  18'd3967,  -18'd10836,  -18'd2275,  18'd5646,  
18'd13813,  -18'd16975,  18'd13802,  18'd13902,  -18'd7948,  -18'd623,  18'd12696,  -18'd15334,  18'd8178,  18'd18869,  18'd1144,  -18'd865,  18'd4300,  18'd3890,  18'd6913,  -18'd1156,  
18'd4653,  18'd2251,  18'd2129,  18'd6254,  18'd4790,  -18'd700,  -18'd7948,  18'd5517,  18'd3013,  -18'd4103,  18'd7363,  18'd12191,  -18'd1015,  -18'd1357,  -18'd5236,  18'd6671,  
-18'd6025,  18'd20716,  18'd5747,  18'd7084,  -18'd1703,  18'd874,  18'd11202,  18'd4276,  -18'd5603,  -18'd5022,  18'd8717,  18'd4324,  18'd6515,  18'd336,  18'd4036,  18'd1863,  
18'd1051,  18'd15523,  18'd16496,  18'd3216,  -18'd8321,  18'd11691,  18'd19545,  18'd4807,  18'd14622,  -18'd7634,  -18'd6796,  -18'd10639,  18'd4926,  -18'd11744,  18'd7137,  18'd7317,  
-18'd592,  18'd6972,  18'd24412,  -18'd9973,  18'd1329,  18'd14731,  18'd8993,  18'd627,  -18'd8890,  18'd8089,  -18'd585,  -18'd14621,  -18'd3250,  -18'd2503,  18'd3672,  -18'd10281,  
18'd8480,  18'd9675,  -18'd1326,  18'd21676,  -18'd4203,  -18'd5954,  -18'd4832,  -18'd15294,  18'd3937,  -18'd7858,  -18'd1371,  18'd14118,  -18'd6330,  18'd15455,  -18'd11229,  18'd24130,  
18'd2268,  18'd13108,  -18'd11050,  18'd12641,  -18'd2143,  -18'd1942,  -18'd17317,  -18'd1488,  18'd15221,  -18'd2721,  -18'd6598,  18'd13125,  -18'd8081,  18'd10193,  -18'd3816,  18'd483,  
-18'd3880,  18'd7758,  18'd7918,  18'd3929,  -18'd2750,  -18'd7349,  18'd3505,  18'd12589,  18'd582,  18'd945,  -18'd2800,  -18'd17291,  18'd3613,  18'd4551,  18'd332,  18'd12800,  
-18'd9696,  18'd21780,  18'd11669,  -18'd7183,  -18'd4430,  18'd5108,  -18'd6200,  18'd17930,  -18'd23627,  -18'd7891,  18'd8976,  -18'd1993,  -18'd8890,  18'd13716,  -18'd1955,  -18'd3546,  

18'd20438,  -18'd1195,  18'd1585,  18'd12471,  18'd1589,  18'd13042,  18'd7993,  -18'd1466,  18'd804,  18'd3826,  18'd11099,  18'd12353,  -18'd5033,  18'd5189,  -18'd4541,  18'd13327,  
18'd2607,  18'd2377,  18'd1266,  18'd23927,  18'd1124,  -18'd4629,  18'd7936,  18'd721,  18'd5883,  -18'd5701,  18'd11490,  -18'd6698,  -18'd12321,  -18'd14884,  18'd17066,  -18'd5109,  
18'd7060,  -18'd119,  18'd17247,  18'd4185,  18'd7962,  -18'd4153,  18'd10416,  18'd12427,  -18'd2987,  -18'd10108,  18'd9385,  -18'd12995,  -18'd12732,  -18'd23961,  18'd13420,  18'd8837,  
-18'd10700,  18'd514,  18'd4874,  18'd2181,  -18'd1564,  -18'd11023,  18'd23431,  18'd10204,  -18'd13344,  -18'd8716,  -18'd11610,  -18'd13800,  -18'd8671,  -18'd7200,  -18'd5,  18'd8053,  
18'd2156,  18'd9584,  18'd11358,  18'd10595,  18'd1458,  18'd7416,  18'd9640,  -18'd6381,  18'd2383,  18'd5841,  -18'd422,  -18'd3279,  -18'd1967,  -18'd9307,  18'd9382,  -18'd4072,  
18'd710,  -18'd3419,  18'd11642,  18'd10535,  18'd1668,  18'd8176,  18'd12107,  -18'd2282,  18'd10449,  18'd10713,  18'd5422,  18'd9651,  18'd3041,  -18'd1750,  18'd4123,  -18'd1932,  
18'd10121,  18'd6904,  18'd5868,  18'd1304,  -18'd7758,  18'd7827,  18'd497,  18'd9931,  18'd5067,  -18'd15547,  18'd4491,  18'd5762,  18'd3395,  -18'd1703,  -18'd11520,  -18'd5235,  
-18'd6119,  18'd5784,  18'd4418,  -18'd2902,  18'd7598,  18'd3732,  -18'd2816,  18'd4711,  -18'd20367,  18'd13234,  -18'd8226,  -18'd2893,  -18'd3925,  18'd6071,  18'd1066,  18'd11414,  
18'd1352,  18'd8344,  18'd5219,  18'd1961,  -18'd3131,  -18'd14804,  -18'd5168,  18'd3929,  -18'd14400,  18'd7197,  18'd3149,  18'd14814,  18'd2977,  18'd14731,  -18'd996,  18'd3751,  
-18'd9422,  -18'd1872,  18'd12545,  -18'd2879,  -18'd7701,  -18'd3439,  18'd12616,  18'd15767,  18'd12857,  18'd9133,  18'd5142,  18'd5125,  -18'd1776,  18'd9099,  -18'd9466,  -18'd1328,  
-18'd8991,  -18'd124,  -18'd368,  -18'd677,  -18'd840,  18'd8080,  -18'd9611,  -18'd12312,  -18'd7040,  -18'd9897,  -18'd3108,  18'd2646,  -18'd239,  18'd2497,  -18'd14660,  -18'd7137,  
-18'd1568,  18'd7501,  -18'd20793,  18'd2363,  18'd6279,  18'd4209,  18'd2551,  18'd1871,  18'd2918,  -18'd10627,  -18'd20542,  -18'd9198,  -18'd7781,  18'd12400,  -18'd11499,  -18'd4993,  
-18'd5650,  18'd9859,  -18'd10688,  18'd15165,  -18'd912,  -18'd17103,  -18'd7098,  18'd13614,  18'd1349,  18'd8439,  -18'd802,  18'd10497,  18'd228,  18'd10680,  18'd10635,  18'd4789,  
-18'd5128,  18'd12746,  18'd4790,  -18'd5577,  18'd1564,  -18'd2382,  -18'd6967,  18'd14051,  -18'd4245,  18'd14544,  18'd9945,  -18'd3700,  -18'd5638,  18'd22108,  18'd1316,  -18'd369,  
-18'd9308,  -18'd559,  18'd3734,  18'd3963,  -18'd4846,  18'd22248,  18'd14098,  -18'd12785,  -18'd7577,  -18'd474,  -18'd7950,  18'd1186,  18'd4069,  18'd21262,  18'd838,  18'd1494,  
18'd12088,  -18'd28722,  -18'd20283,  -18'd2283,  18'd5380,  18'd29325,  -18'd2417,  -18'd17338,  18'd12115,  -18'd8042,  -18'd13244,  18'd9059,  18'd173,  18'd17015,  18'd3569,  18'd1459,  

18'd2464,  -18'd29520,  -18'd11103,  18'd3298,  -18'd4735,  18'd6081,  18'd11230,  -18'd6689,  18'd3152,  18'd19687,  -18'd16219,  -18'd8142,  18'd3712,  -18'd2963,  -18'd12783,  -18'd25135,  
18'd19101,  -18'd26795,  18'd2240,  18'd7618,  18'd4633,  -18'd4036,  18'd6852,  -18'd11194,  -18'd880,  18'd18364,  18'd3643,  -18'd1476,  18'd2229,  18'd6846,  -18'd11244,  -18'd6476,  
18'd9931,  -18'd3959,  -18'd13283,  -18'd16037,  18'd6057,  18'd7528,  18'd26307,  18'd2061,  18'd15603,  -18'd4349,  18'd3516,  18'd22644,  -18'd5048,  -18'd1933,  18'd2867,  -18'd22654,  
18'd14161,  18'd343,  18'd22668,  -18'd19301,  18'd4818,  18'd9584,  -18'd789,  18'd412,  18'd12857,  -18'd19693,  -18'd8589,  18'd20645,  -18'd1647,  18'd269,  -18'd10358,  -18'd7547,  
18'd21821,  -18'd24212,  18'd3956,  18'd13170,  18'd5456,  18'd13719,  18'd4740,  18'd80,  18'd2764,  18'd5529,  -18'd5042,  18'd7247,  18'd9438,  18'd1811,  -18'd1908,  -18'd8956,  
18'd3589,  -18'd6165,  -18'd8717,  18'd2273,  18'd6551,  18'd6928,  18'd5736,  -18'd10981,  18'd3152,  18'd1303,  18'd2757,  18'd4852,  18'd5778,  -18'd9538,  -18'd12156,  18'd1516,  
18'd11812,  -18'd3990,  -18'd13377,  -18'd8991,  18'd4263,  -18'd11113,  18'd4526,  18'd7481,  -18'd6134,  -18'd5742,  -18'd9285,  18'd8307,  -18'd196,  18'd10549,  -18'd4773,  18'd12334,  
-18'd13989,  18'd4909,  18'd9029,  -18'd13062,  18'd4389,  -18'd5997,  -18'd11580,  18'd20964,  18'd1982,  -18'd3907,  18'd8001,  18'd3388,  -18'd1509,  18'd2473,  18'd2894,  18'd10872,  
18'd3192,  -18'd6488,  18'd3544,  -18'd14156,  18'd4036,  18'd5036,  18'd521,  -18'd1736,  18'd2608,  -18'd18482,  18'd2475,  18'd8315,  -18'd5866,  -18'd2532,  -18'd1604,  18'd2277,  
18'd0,  18'd12190,  -18'd10533,  18'd5480,  18'd8579,  18'd256,  18'd7757,  -18'd4537,  -18'd639,  -18'd6371,  18'd2775,  -18'd1284,  18'd8629,  18'd7542,  18'd9781,  18'd9046,  
18'd4148,  18'd8923,  -18'd13034,  18'd3576,  -18'd7706,  18'd7268,  18'd3534,  -18'd186,  -18'd366,  -18'd4677,  18'd6119,  18'd9442,  -18'd5544,  -18'd9309,  18'd3959,  -18'd5327,  
-18'd954,  18'd3601,  18'd8673,  -18'd5316,  -18'd7430,  -18'd11532,  -18'd6559,  18'd12198,  -18'd5602,  18'd8444,  18'd18806,  18'd15436,  -18'd6579,  -18'd359,  -18'd10595,  18'd6901,  
18'd15682,  18'd9104,  18'd5598,  18'd3005,  18'd2225,  18'd14936,  18'd3277,  18'd10702,  18'd13063,  -18'd6784,  18'd17516,  -18'd12410,  18'd7925,  -18'd4145,  -18'd32,  18'd10500,  
18'd1086,  -18'd13376,  18'd16963,  18'd7997,  18'd5330,  18'd1783,  18'd11862,  -18'd4463,  18'd4021,  -18'd18295,  18'd4842,  -18'd1130,  -18'd6758,  -18'd8193,  18'd10867,  -18'd6225,  
-18'd4508,  -18'd18432,  18'd22978,  18'd4915,  -18'd3986,  -18'd11497,  -18'd1273,  18'd13242,  18'd6386,  18'd21034,  18'd8171,  -18'd2876,  -18'd4769,  -18'd17140,  18'd13128,  -18'd5760,  
-18'd6860,  18'd17906,  18'd1284,  18'd4924,  18'd5183,  -18'd12210,  18'd6559,  18'd10904,  -18'd16676,  18'd15167,  18'd10445,  18'd7128,  -18'd656,  18'd535,  18'd16626,  18'd740,  

-18'd5074,  -18'd10457,  18'd4497,  18'd7461,  18'd1069,  -18'd3806,  -18'd7055,  -18'd3768,  18'd4215,  18'd14664,  -18'd9049,  18'd2028,  -18'd5744,  18'd3806,  18'd6781,  18'd1452,  
18'd95,  -18'd6272,  -18'd7332,  18'd6038,  18'd6945,  -18'd17706,  18'd559,  -18'd2171,  -18'd23849,  -18'd15014,  -18'd10329,  -18'd6163,  18'd6260,  18'd4434,  -18'd8841,  -18'd6673,  
-18'd11649,  -18'd9462,  18'd3163,  18'd38,  -18'd4367,  18'd6801,  -18'd6467,  18'd1768,  -18'd9645,  -18'd13178,  -18'd8757,  -18'd4802,  18'd4117,  -18'd259,  18'd10130,  -18'd15895,  
-18'd10655,  -18'd4311,  18'd12911,  -18'd5150,  -18'd6317,  -18'd10447,  18'd836,  18'd1598,  -18'd16880,  -18'd4133,  -18'd8005,  -18'd13044,  18'd5682,  -18'd7695,  18'd204,  -18'd11147,  
-18'd3332,  -18'd8131,  -18'd8958,  18'd7357,  -18'd8193,  -18'd951,  -18'd5234,  -18'd3348,  -18'd6416,  18'd8149,  18'd2226,  18'd6470,  -18'd9502,  18'd6384,  18'd10421,  -18'd7368,  
18'd802,  -18'd8745,  -18'd1452,  18'd18477,  18'd4367,  -18'd7625,  -18'd13623,  -18'd5590,  -18'd10622,  -18'd4691,  18'd6391,  18'd6181,  18'd7576,  18'd1660,  18'd2337,  -18'd6742,  
-18'd911,  18'd4558,  -18'd1612,  -18'd5653,  18'd236,  -18'd937,  18'd1794,  -18'd1948,  18'd19,  -18'd11533,  18'd5938,  18'd9858,  18'd4337,  -18'd6999,  18'd929,  -18'd4292,  
18'd11997,  18'd10131,  18'd1869,  -18'd7127,  -18'd1684,  -18'd7072,  18'd7818,  18'd10237,  -18'd6441,  18'd271,  18'd3498,  -18'd8466,  -18'd8973,  18'd6194,  18'd5846,  -18'd6600,  
-18'd3429,  -18'd1713,  -18'd16185,  -18'd9601,  -18'd4203,  -18'd5063,  -18'd8161,  -18'd4889,  -18'd7849,  -18'd4587,  18'd11067,  -18'd5917,  18'd1331,  18'd3215,  -18'd2211,  -18'd12362,  
-18'd13431,  18'd8090,  -18'd6520,  18'd3185,  -18'd3226,  18'd1248,  -18'd5873,  18'd10064,  -18'd9443,  -18'd6123,  18'd10401,  -18'd3016,  18'd5712,  18'd6790,  18'd3594,  -18'd1656,  
-18'd3334,  18'd969,  -18'd2631,  18'd4825,  -18'd7069,  -18'd1869,  -18'd4909,  -18'd6175,  -18'd3099,  -18'd3298,  -18'd14479,  18'd6113,  -18'd5059,  18'd4099,  -18'd6590,  -18'd2834,  
18'd2838,  18'd12868,  -18'd6523,  -18'd6638,  -18'd694,  -18'd9439,  -18'd17192,  -18'd3697,  -18'd4428,  18'd1251,  -18'd11510,  18'd13540,  -18'd7599,  18'd6289,  -18'd20482,  18'd13648,  
18'd5828,  -18'd11742,  -18'd11917,  -18'd7801,  -18'd3880,  18'd1258,  18'd9306,  -18'd13031,  -18'd6595,  18'd1849,  18'd7636,  18'd7784,  -18'd2135,  18'd417,  18'd1726,  18'd448,  
18'd7052,  18'd319,  18'd3160,  -18'd2359,  18'd7099,  18'd1287,  -18'd14474,  -18'd5875,  -18'd10428,  -18'd8895,  -18'd9593,  -18'd6937,  18'd2854,  18'd3469,  18'd3199,  -18'd10267,  
18'd4576,  -18'd13039,  -18'd9635,  -18'd8678,  -18'd6943,  18'd14113,  -18'd13987,  -18'd9530,  -18'd6340,  18'd1338,  -18'd1368,  18'd7546,  18'd3178,  -18'd3366,  18'd4154,  -18'd1173,  
-18'd3257,  -18'd5380,  -18'd4362,  18'd6833,  -18'd697,  -18'd2774,  -18'd7185,  18'd7106,  18'd2697,  18'd10179,  -18'd7228,  -18'd2413,  -18'd5472,  18'd8220,  -18'd3016,  18'd12071,  

18'd7468,  -18'd8447,  -18'd8591,  -18'd3612,  18'd7829,  18'd444,  18'd6874,  -18'd6638,  -18'd7307,  -18'd5406,  18'd7334,  18'd6186,  18'd6537,  -18'd6572,  18'd3881,  18'd3033,  
-18'd6951,  18'd2125,  -18'd233,  18'd6579,  -18'd4134,  -18'd3048,  18'd5522,  18'd4882,  -18'd10275,  -18'd976,  -18'd8592,  -18'd2946,  -18'd7207,  -18'd3487,  -18'd3680,  -18'd8103,  
-18'd4124,  -18'd269,  18'd8514,  18'd6456,  -18'd6274,  -18'd1977,  18'd973,  -18'd8460,  -18'd3520,  -18'd1248,  -18'd4513,  -18'd9421,  18'd3703,  18'd5542,  -18'd3579,  -18'd5715,  
18'd5864,  -18'd4959,  18'd7447,  18'd4527,  18'd1314,  18'd7708,  18'd1240,  -18'd4123,  -18'd1332,  -18'd9046,  18'd3243,  -18'd1317,  18'd4431,  -18'd4355,  18'd3040,  -18'd9009,  
-18'd1508,  -18'd3410,  -18'd11264,  -18'd1713,  18'd2590,  18'd5160,  18'd2619,  -18'd8994,  18'd4233,  18'd6373,  -18'd6468,  -18'd2138,  -18'd4279,  18'd5279,  18'd4399,  -18'd1897,  
18'd5243,  -18'd6606,  -18'd6744,  18'd4319,  18'd5037,  -18'd2925,  -18'd1252,  18'd2896,  -18'd8602,  -18'd8500,  18'd6623,  -18'd3529,  -18'd5228,  18'd3825,  18'd5503,  18'd4356,  
-18'd3790,  -18'd4855,  -18'd6081,  -18'd4499,  18'd4467,  -18'd9322,  -18'd9274,  18'd6911,  18'd2849,  -18'd1190,  18'd877,  -18'd5132,  -18'd2941,  -18'd8959,  -18'd9945,  18'd2723,  
18'd2542,  -18'd4296,  -18'd4216,  -18'd4874,  -18'd7122,  -18'd5106,  -18'd2081,  18'd5578,  -18'd9536,  -18'd11428,  18'd1311,  -18'd4908,  -18'd8265,  18'd1286,  -18'd9200,  18'd6807,  
-18'd7694,  -18'd257,  -18'd6369,  -18'd401,  18'd1913,  18'd5950,  -18'd739,  -18'd5614,  -18'd6948,  18'd6935,  -18'd344,  -18'd3697,  -18'd3169,  18'd167,  -18'd8936,  -18'd4610,  
-18'd3189,  -18'd8701,  18'd4445,  -18'd6581,  18'd1083,  18'd7841,  18'd1536,  18'd3480,  18'd520,  -18'd5540,  -18'd6430,  -18'd8358,  -18'd7036,  -18'd7080,  -18'd8367,  -18'd9387,  
-18'd3797,  18'd0,  18'd5166,  -18'd9285,  -18'd6054,  -18'd7149,  18'd4722,  18'd6813,  -18'd7980,  -18'd806,  -18'd2862,  -18'd3085,  18'd8529,  -18'd6710,  -18'd6871,  18'd6825,  
18'd1347,  -18'd3031,  -18'd745,  -18'd10426,  18'd458,  18'd8460,  18'd4108,  18'd1533,  -18'd3549,  -18'd10368,  -18'd1445,  -18'd7686,  -18'd1563,  -18'd3081,  18'd1202,  -18'd1620,  
18'd3695,  -18'd8777,  -18'd63,  18'd6940,  18'd1869,  -18'd7128,  -18'd3889,  -18'd9572,  -18'd10729,  -18'd1482,  -18'd2369,  18'd2492,  -18'd6805,  -18'd5510,  -18'd4850,  18'd5611,  
18'd1,  18'd1216,  -18'd5439,  -18'd11889,  18'd7238,  -18'd1332,  -18'd9048,  18'd2279,  -18'd6559,  18'd1823,  18'd5772,  -18'd6884,  18'd5499,  -18'd468,  18'd729,  -18'd9960,  
18'd4069,  -18'd9180,  18'd4120,  18'd6468,  18'd4950,  18'd3311,  -18'd9879,  -18'd2980,  18'd4654,  -18'd3435,  -18'd6775,  -18'd6631,  18'd3085,  18'd6799,  18'd1776,  18'd5641,  
-18'd7736,  18'd1966,  -18'd7495,  -18'd3385,  18'd6409,  -18'd8588,  -18'd7205,  -18'd5917,  -18'd761,  18'd6705,  18'd6874,  -18'd1634,  18'd3789,  18'd3103,  18'd2844,  -18'd1527,  

-18'd9152,  -18'd2833,  18'd10052,  18'd7531,  18'd127,  18'd6275,  -18'd3459,  -18'd451,  18'd15903,  -18'd6236,  18'd8599,  -18'd4179,  -18'd5289,  18'd2478,  18'd10535,  18'd28878,  
-18'd4069,  18'd16597,  18'd5124,  18'd11179,  -18'd1595,  -18'd2399,  18'd692,  18'd18740,  -18'd6488,  18'd4258,  18'd8209,  18'd7722,  18'd1691,  -18'd7551,  18'd3309,  -18'd441,  
-18'd12340,  18'd13133,  -18'd4422,  18'd13165,  18'd1388,  -18'd1132,  18'd15559,  18'd10904,  18'd6884,  -18'd10996,  18'd12895,  -18'd12240,  18'd7642,  -18'd12555,  18'd14114,  -18'd5824,  
-18'd19586,  18'd14849,  -18'd20493,  18'd2147,  -18'd5808,  -18'd9791,  18'd4494,  18'd15081,  -18'd25496,  18'd14134,  18'd7869,  18'd2102,  18'd7479,  -18'd4773,  18'd3099,  18'd4454,  
18'd16071,  18'd15220,  18'd3547,  -18'd14542,  18'd2129,  18'd6571,  -18'd4302,  -18'd500,  18'd15448,  -18'd16191,  -18'd341,  18'd6884,  18'd10100,  18'd9617,  -18'd6523,  18'd15788,  
18'd24821,  -18'd12268,  18'd4824,  18'd21731,  -18'd5491,  -18'd2698,  -18'd6585,  -18'd5744,  18'd11840,  -18'd5268,  -18'd11970,  -18'd1584,  18'd3954,  -18'd514,  -18'd12011,  -18'd62,  
18'd3071,  -18'd18029,  -18'd11403,  18'd4049,  18'd2530,  -18'd1694,  18'd15697,  18'd16579,  18'd3212,  18'd10295,  -18'd17903,  18'd13674,  -18'd5548,  -18'd5035,  18'd8682,  -18'd18630,  
18'd3727,  -18'd7355,  -18'd3278,  -18'd4175,  -18'd8789,  18'd9408,  18'd18031,  -18'd11576,  18'd5345,  -18'd2317,  18'd25413,  -18'd7257,  -18'd3611,  -18'd17442,  18'd16621,  -18'd10061,  
18'd26015,  -18'd6998,  18'd6812,  18'd7866,  -18'd6692,  18'd2174,  18'd2486,  -18'd13515,  18'd6860,  -18'd3437,  18'd1843,  -18'd4682,  -18'd470,  18'd2716,  18'd1761,  -18'd11441,  
18'd12472,  -18'd16732,  18'd9053,  -18'd13988,  -18'd8305,  18'd6246,  18'd6311,  -18'd7672,  18'd6334,  18'd3159,  18'd9317,  -18'd1974,  18'd10509,  -18'd3393,  18'd4755,  -18'd2287,  
18'd551,  -18'd1968,  -18'd16434,  18'd3755,  18'd3785,  -18'd14256,  -18'd10210,  18'd1220,  -18'd12017,  18'd9965,  -18'd21536,  18'd4092,  -18'd6503,  -18'd9814,  -18'd4826,  18'd2855,  
18'd7752,  -18'd10989,  18'd8549,  -18'd771,  -18'd9294,  18'd6712,  18'd13452,  18'd9529,  -18'd17870,  -18'd21843,  18'd8934,  -18'd7772,  18'd1092,  -18'd15238,  18'd2665,  -18'd14306,  
18'd15659,  -18'd11005,  18'd3374,  -18'd13249,  18'd7731,  -18'd7226,  -18'd2690,  -18'd12527,  18'd6052,  -18'd12461,  -18'd5225,  -18'd2393,  18'd5120,  -18'd1228,  -18'd11407,  -18'd5866,  
-18'd14941,  18'd384,  18'd15375,  -18'd2209,  -18'd5439,  18'd15154,  -18'd4330,  18'd21007,  18'd11812,  18'd4264,  18'd2231,  18'd8604,  18'd9776,  18'd2760,  -18'd12707,  18'd15058,  
-18'd1656,  18'd13262,  18'd3377,  18'd10506,  18'd5321,  -18'd15531,  -18'd8083,  -18'd3246,  -18'd1591,  -18'd67,  -18'd7968,  -18'd5409,  18'd714,  -18'd2064,  -18'd13782,  18'd2195,  
18'd9735,  18'd3340,  18'd9877,  -18'd644,  -18'd7707,  18'd8642,  18'd5032,  -18'd1329,  -18'd15744,  -18'd14456,  -18'd8812,  18'd3834,  -18'd312,  18'd751,  -18'd3233,  -18'd3377,  

18'd28180,  18'd19885,  18'd9758,  18'd23584,  18'd6400,  -18'd3574,  18'd10640,  -18'd263,  18'd7221,  -18'd19438,  18'd13054,  -18'd6707,  18'd2257,  18'd3180,  -18'd369,  18'd23683,  
-18'd6273,  18'd6762,  -18'd1023,  -18'd16186,  18'd3,  -18'd14032,  -18'd2134,  18'd2246,  -18'd11176,  -18'd14693,  -18'd21180,  -18'd28589,  18'd5284,  -18'd13626,  18'd23576,  18'd5105,  
18'd582,  18'd317,  18'd28081,  -18'd9415,  -18'd7980,  18'd27376,  18'd24810,  18'd15754,  -18'd3780,  18'd1078,  18'd1381,  -18'd3681,  18'd2288,  -18'd2445,  18'd3936,  18'd10626,  
-18'd20088,  18'd5574,  18'd8840,  -18'd6048,  -18'd4974,  18'd14594,  -18'd411,  -18'd6158,  18'd12554,  18'd14263,  -18'd10377,  18'd205,  18'd6252,  18'd4560,  -18'd2290,  18'd16958,  
18'd5917,  18'd3656,  18'd39,  18'd22188,  -18'd7325,  18'd1212,  -18'd2660,  18'd1194,  18'd16551,  -18'd12200,  -18'd4472,  18'd4174,  -18'd71,  -18'd2244,  18'd3574,  18'd6948,  
18'd13716,  -18'd12071,  -18'd9106,  -18'd3833,  -18'd4539,  -18'd9009,  18'd3595,  18'd2617,  -18'd11992,  -18'd8020,  -18'd3206,  18'd3473,  18'd5042,  18'd962,  18'd3521,  -18'd9011,  
18'd2775,  18'd6677,  18'd14155,  -18'd14174,  -18'd8085,  18'd10356,  18'd19002,  18'd19198,  -18'd1690,  18'd8095,  18'd3110,  18'd7534,  -18'd686,  -18'd7176,  18'd16932,  -18'd9154,  
18'd3156,  18'd18903,  -18'd2062,  18'd2536,  18'd6519,  18'd22750,  18'd14461,  18'd1676,  18'd5774,  -18'd13690,  18'd8872,  -18'd5617,  -18'd3381,  18'd8166,  18'd9149,  18'd2270,  
-18'd8425,  18'd10741,  -18'd3165,  18'd17024,  -18'd5329,  18'd11817,  18'd996,  18'd11503,  -18'd1309,  -18'd9969,  -18'd7358,  -18'd8421,  -18'd5853,  18'd7119,  -18'd7593,  18'd5662,  
18'd9990,  -18'd11970,  -18'd7597,  18'd15849,  18'd3368,  18'd3563,  -18'd9121,  18'd1469,  -18'd5861,  18'd12000,  -18'd15105,  -18'd8870,  -18'd4306,  -18'd8935,  -18'd19665,  18'd4279,  
18'd1242,  -18'd6747,  -18'd17026,  -18'd1276,  -18'd6497,  -18'd7060,  -18'd8465,  -18'd7152,  -18'd13387,  -18'd10705,  -18'd7277,  -18'd8643,  -18'd6612,  -18'd8070,  18'd3505,  -18'd7640,  
18'd8272,  18'd22207,  -18'd3362,  -18'd668,  -18'd7821,  18'd16188,  -18'd5396,  18'd14174,  18'd16975,  -18'd12782,  18'd220,  -18'd3370,  18'd7539,  18'd12403,  18'd7729,  18'd8524,  
18'd10634,  18'd25948,  -18'd8816,  18'd16227,  18'd4731,  18'd11134,  -18'd2779,  18'd23372,  -18'd1402,  -18'd267,  -18'd1689,  18'd17844,  18'd4449,  18'd13976,  18'd6247,  18'd8380,  
-18'd11566,  18'd4274,  18'd1541,  18'd16785,  18'd276,  -18'd2715,  -18'd2356,  18'd2569,  -18'd898,  18'd5089,  18'd7922,  -18'd695,  -18'd6608,  18'd15627,  -18'd11975,  18'd9080,  
18'd5081,  18'd9666,  -18'd15407,  18'd5911,  18'd6243,  -18'd15497,  -18'd9309,  -18'd11053,  -18'd20272,  -18'd197,  -18'd3286,  -18'd9810,  -18'd4190,  -18'd4976,  18'd2695,  -18'd691,  
-18'd2402,  18'd8190,  -18'd6578,  -18'd2564,  18'd2946,  18'd24080,  -18'd8545,  -18'd708,  -18'd5864,  -18'd19255,  -18'd10861,  -18'd5189,  -18'd6931,  18'd5907,  18'd11944,  18'd777,  

18'd567,  -18'd9631,  18'd17268,  -18'd4203,  18'd7343,  18'd18272,  18'd4446,  -18'd4031,  18'd7821,  18'd5545,  18'd1601,  18'd6809,  -18'd7739,  18'd2984,  -18'd521,  -18'd4522,  
18'd10681,  18'd804,  18'd1371,  18'd20148,  -18'd5218,  18'd9393,  -18'd5623,  -18'd18579,  18'd11866,  -18'd8379,  -18'd3405,  18'd7550,  18'd5725,  18'd11470,  18'd3542,  -18'd23475,  
18'd13861,  -18'd15434,  -18'd17941,  18'd20442,  -18'd6390,  -18'd10624,  -18'd14017,  -18'd11164,  18'd9525,  18'd991,  -18'd13956,  18'd4509,  18'd4842,  -18'd19821,  -18'd14348,  -18'd1544,  
18'd8508,  -18'd21876,  -18'd17918,  -18'd20594,  18'd6502,  -18'd11253,  18'd14605,  18'd23107,  18'd8522,  -18'd12580,  -18'd17534,  -18'd18200,  18'd2554,  -18'd4980,  -18'd8169,  -18'd28543,  
-18'd8050,  18'd20277,  18'd16471,  18'd2735,  -18'd3564,  18'd5523,  -18'd5339,  18'd6315,  18'd8127,  -18'd30530,  18'd5390,  -18'd70,  -18'd3231,  -18'd4297,  -18'd2366,  18'd7186,  
18'd5085,  18'd5809,  18'd1096,  -18'd4205,  18'd6612,  18'd5652,  18'd10978,  18'd1813,  18'd6775,  18'd1397,  18'd7626,  -18'd8471,  18'd1949,  18'd6157,  -18'd2669,  18'd14932,  
-18'd1898,  18'd12185,  -18'd24593,  18'd12469,  -18'd3542,  -18'd20600,  -18'd6013,  -18'd8398,  -18'd6987,  18'd3037,  -18'd20729,  -18'd10245,  18'd15,  18'd1823,  -18'd2606,  18'd7109,  
18'd12531,  -18'd21348,  -18'd17782,  18'd499,  -18'd3168,  18'd9113,  18'd11482,  18'd1338,  -18'd37814,  -18'd18643,  -18'd11324,  -18'd13884,  18'd7902,  -18'd1414,  -18'd4343,  -18'd4283,  
-18'd9362,  18'd18459,  18'd5420,  18'd17156,  18'd7610,  18'd9764,  -18'd8649,  18'd8800,  18'd7558,  18'd604,  18'd2520,  18'd13368,  -18'd2581,  18'd3579,  -18'd10940,  18'd18041,  
18'd3140,  18'd7092,  18'd9282,  18'd5667,  18'd6129,  18'd7077,  -18'd17217,  -18'd9851,  18'd4620,  -18'd1839,  -18'd11842,  18'd11615,  -18'd4996,  18'd20472,  18'd166,  18'd10199,  
-18'd167,  -18'd527,  -18'd19776,  18'd10995,  18'd1267,  18'd992,  18'd1587,  -18'd24387,  -18'd10120,  -18'd12756,  18'd6608,  -18'd12429,  18'd4196,  -18'd3030,  18'd8102,  18'd3235,  
18'd6604,  -18'd44770,  18'd502,  18'd6228,  -18'd1227,  18'd1554,  18'd13374,  -18'd7724,  -18'd27533,  -18'd16134,  18'd16551,  -18'd672,  -18'd7148,  -18'd11698,  18'd6540,  -18'd17684,  
-18'd2683,  18'd4804,  18'd7538,  18'd9636,  -18'd7470,  18'd12594,  -18'd6034,  18'd5741,  18'd9495,  18'd3661,  18'd641,  -18'd692,  18'd1750,  18'd10673,  -18'd4399,  18'd5683,  
18'd9742,  18'd2073,  -18'd6872,  18'd10721,  18'd400,  18'd15755,  -18'd19286,  -18'd12908,  18'd1213,  18'd10189,  -18'd3562,  18'd11195,  -18'd7892,  18'd7697,  -18'd6213,  18'd13684,  
18'd1780,  -18'd11289,  -18'd8059,  18'd12130,  -18'd3870,  18'd5936,  18'd8166,  -18'd10947,  18'd7906,  18'd2206,  -18'd3696,  -18'd2414,  18'd5908,  -18'd15021,  18'd16217,  18'd12265,  
18'd4246,  -18'd3921,  18'd16529,  -18'd8766,  -18'd5326,  -18'd326,  18'd25883,  -18'd5126,  -18'd1780,  -18'd24966,  18'd9302,  -18'd20040,  18'd4046,  -18'd28042,  18'd6868,  18'd942,  

18'd3716,  -18'd15613,  18'd1114,  -18'd22334,  18'd3377,  18'd3324,  18'd12065,  -18'd7896,  18'd14024,  18'd13092,  18'd992,  18'd9727,  18'd5161,  -18'd10519,  -18'd2624,  -18'd15539,  
18'd17808,  -18'd8808,  -18'd4332,  -18'd7211,  -18'd1926,  18'd14762,  18'd10997,  18'd1028,  18'd22931,  18'd24500,  18'd10443,  18'd29040,  18'd1673,  18'd18546,  -18'd10229,  -18'd5358,  
18'd5754,  -18'd3480,  18'd757,  18'd11195,  -18'd589,  18'd7185,  18'd13846,  -18'd15793,  18'd20137,  18'd15206,  -18'd10208,  18'd20328,  18'd4753,  18'd12025,  -18'd7695,  -18'd8633,  
18'd10067,  -18'd3633,  18'd9209,  18'd16380,  18'd2823,  -18'd9979,  -18'd9164,  18'd6006,  18'd20232,  -18'd5038,  -18'd12637,  18'd17039,  18'd7060,  -18'd5311,  -18'd11176,  18'd10372,  
-18'd3332,  -18'd2194,  -18'd10202,  18'd977,  18'd66,  18'd5488,  18'd8550,  18'd10082,  18'd12633,  -18'd982,  18'd11341,  -18'd11757,  -18'd95,  18'd3561,  -18'd398,  18'd2927,  
-18'd3072,  -18'd3761,  -18'd657,  18'd5512,  -18'd4862,  18'd6574,  18'd6728,  -18'd12527,  18'd9651,  -18'd8579,  18'd868,  18'd1404,  18'd5298,  -18'd188,  -18'd5687,  18'd4470,  
18'd7532,  -18'd5041,  -18'd6412,  -18'd6814,  -18'd7142,  -18'd556,  18'd884,  -18'd17435,  -18'd16062,  18'd18694,  -18'd15633,  18'd1113,  -18'd767,  18'd1222,  18'd8752,  -18'd8882,  
-18'd6862,  -18'd11175,  -18'd12723,  18'd8569,  18'd3381,  -18'd11152,  -18'd9878,  18'd1417,  18'd15387,  18'd2112,  -18'd559,  18'd292,  -18'd3855,  18'd3735,  18'd8407,  -18'd18269,  
18'd10287,  -18'd3286,  18'd3617,  18'd21946,  -18'd1968,  18'd11581,  18'd12895,  18'd11167,  18'd8458,  -18'd160,  18'd7136,  -18'd3883,  18'd12775,  -18'd14972,  18'd13621,  18'd2089,  
18'd856,  18'd866,  -18'd491,  -18'd9823,  18'd5682,  -18'd4795,  18'd6320,  -18'd9953,  -18'd1929,  18'd3461,  18'd54,  -18'd12879,  18'd12598,  -18'd10956,  -18'd562,  18'd4546,  
18'd8827,  18'd1496,  -18'd6413,  -18'd3950,  -18'd2085,  -18'd429,  18'd1803,  18'd1121,  -18'd10566,  18'd1651,  -18'd7150,  -18'd15471,  18'd2089,  -18'd2795,  -18'd893,  18'd2391,  
-18'd6914,  18'd2537,  -18'd10521,  18'd3244,  -18'd1171,  -18'd10626,  18'd1973,  -18'd810,  -18'd3917,  -18'd14124,  -18'd1666,  18'd965,  -18'd1457,  -18'd1526,  18'd9123,  -18'd10848,  
18'd27995,  18'd11720,  18'd7550,  18'd9460,  -18'd6693,  18'd7167,  -18'd6783,  18'd15649,  18'd3273,  18'd7030,  18'd4,  18'd14231,  18'd10645,  -18'd7106,  -18'd6437,  -18'd4937,  
-18'd3062,  -18'd19560,  18'd9058,  -18'd9449,  18'd1982,  18'd12612,  18'd14871,  18'd2889,  18'd9292,  -18'd2457,  18'd12763,  18'd3692,  -18'd4289,  -18'd19821,  -18'd1495,  18'd3205,  
18'd16585,  -18'd22204,  18'd8033,  -18'd1629,  18'd461,  18'd5493,  18'd10303,  18'd8542,  18'd13931,  18'd1570,  18'd5342,  18'd8708,  -18'd4395,  -18'd9527,  18'd5298,  -18'd16837,  
18'd15562,  -18'd730,  18'd11092,  -18'd3400,  -18'd2236,  18'd2496,  18'd6989,  18'd10431,  18'd15282,  -18'd5529,  18'd7406,  18'd770,  18'd680,  18'd5335,  18'd4020,  -18'd12388,  

-18'd4150,  -18'd5349,  18'd5956,  -18'd7486,  -18'd2391,  18'd1197,  18'd774,  -18'd4910,  -18'd2553,  -18'd7928,  -18'd7090,  -18'd1376,  18'd1620,  -18'd7703,  -18'd4588,  -18'd4694,  
18'd1704,  18'd4316,  18'd5511,  18'd3123,  -18'd2279,  -18'd8989,  18'd1540,  -18'd8340,  -18'd6312,  -18'd10410,  18'd1540,  18'd4934,  -18'd7895,  18'd145,  -18'd3676,  18'd3805,  
-18'd8495,  -18'd11500,  -18'd9915,  18'd1713,  -18'd722,  -18'd6893,  18'd5617,  -18'd5545,  18'd1007,  -18'd2818,  18'd2006,  -18'd8592,  -18'd3107,  -18'd8050,  18'd6093,  -18'd7473,  
-18'd9340,  18'd7626,  -18'd5649,  -18'd1066,  -18'd7713,  -18'd7293,  -18'd4219,  18'd6018,  -18'd3452,  -18'd9752,  18'd1289,  -18'd6011,  -18'd100,  -18'd5986,  -18'd7553,  -18'd5961,  
-18'd5804,  -18'd10613,  18'd5936,  -18'd5683,  -18'd3786,  18'd4528,  18'd5981,  -18'd8385,  -18'd3938,  -18'd8342,  18'd5843,  -18'd11316,  18'd8575,  18'd6154,  18'd863,  -18'd3940,  
18'd8132,  -18'd188,  18'd3565,  18'd5326,  -18'd6365,  -18'd8319,  -18'd1299,  -18'd9038,  18'd3513,  18'd2370,  -18'd1303,  -18'd7854,  18'd1192,  -18'd10489,  -18'd2053,  -18'd2662,  
-18'd1603,  18'd5173,  18'd5929,  -18'd2332,  -18'd4771,  18'd829,  18'd6576,  -18'd7037,  -18'd3868,  -18'd1327,  -18'd7047,  18'd3757,  -18'd1294,  18'd2570,  18'd3203,  18'd2408,  
-18'd724,  18'd4944,  18'd2680,  18'd2924,  -18'd522,  18'd6782,  -18'd8759,  -18'd10577,  -18'd2276,  18'd2172,  18'd6775,  -18'd2717,  18'd1206,  18'd2639,  18'd1523,  18'd3199,  
-18'd5672,  -18'd4792,  -18'd2683,  -18'd6751,  18'd591,  -18'd2416,  18'd1248,  18'd3518,  -18'd8726,  -18'd10316,  -18'd3726,  -18'd8676,  18'd5337,  -18'd8043,  18'd5556,  18'd571,  
-18'd8966,  -18'd6545,  -18'd1255,  -18'd9037,  -18'd5707,  -18'd2170,  -18'd3308,  18'd1594,  -18'd5985,  -18'd3272,  18'd7043,  -18'd8526,  18'd219,  -18'd7597,  18'd1177,  -18'd7587,  
-18'd3483,  18'd1089,  18'd4224,  -18'd8031,  -18'd8497,  -18'd9834,  -18'd10476,  -18'd8750,  -18'd6277,  -18'd5681,  -18'd4683,  18'd4257,  -18'd3792,  -18'd8440,  18'd3344,  -18'd7572,  
18'd6731,  -18'd9161,  18'd6824,  -18'd8321,  18'd8001,  18'd260,  -18'd5583,  18'd6078,  -18'd5526,  18'd876,  -18'd3625,  -18'd8040,  18'd3429,  -18'd6423,  -18'd8641,  -18'd8339,  
-18'd10368,  18'd3238,  18'd6555,  -18'd6210,  -18'd195,  18'd1992,  18'd2310,  -18'd4806,  -18'd8965,  18'd2043,  -18'd108,  18'd3488,  18'd2199,  18'd4247,  -18'd4975,  18'd7283,  
18'd1000,  -18'd2968,  -18'd6609,  18'd545,  -18'd7400,  -18'd10197,  18'd4453,  -18'd4125,  18'd3627,  18'd4507,  18'd6455,  18'd3483,  18'd3369,  18'd16,  -18'd2079,  -18'd8982,  
18'd1549,  -18'd11381,  -18'd6406,  -18'd5477,  18'd1646,  18'd5939,  18'd4927,  18'd5179,  -18'd2163,  -18'd12252,  18'd4074,  18'd4277,  18'd1866,  -18'd10011,  -18'd7461,  -18'd9472,  
18'd1596,  -18'd8955,  18'd2387,  -18'd3772,  18'd793,  18'd4440,  -18'd1313,  -18'd3232,  -18'd7753,  -18'd6858,  18'd1211,  -18'd3492,  -18'd2963,  18'd234,  18'd252,  18'd4604,  

18'd1577,  -18'd8698,  -18'd6153,  -18'd1480,  18'd2820,  18'd6215,  -18'd4428,  -18'd7410,  -18'd4886,  18'd3803,  -18'd9717,  -18'd3526,  -18'd3526,  -18'd7775,  18'd4114,  -18'd1169,  
-18'd4385,  -18'd5389,  -18'd151,  18'd4826,  18'd288,  -18'd3486,  18'd1869,  18'd6116,  18'd2716,  -18'd2387,  -18'd6272,  -18'd2718,  -18'd2816,  18'd3210,  -18'd9941,  18'd6646,  
18'd565,  -18'd3348,  -18'd9330,  -18'd6342,  18'd5060,  -18'd7447,  18'd5905,  -18'd2574,  -18'd3962,  -18'd10051,  -18'd829,  18'd7532,  -18'd2729,  18'd5284,  -18'd3041,  18'd7574,  
-18'd1338,  -18'd1159,  18'd6204,  -18'd5110,  -18'd3124,  18'd5708,  18'd7531,  18'd3248,  18'd503,  -18'd2726,  18'd2101,  -18'd8932,  -18'd4908,  -18'd3727,  18'd1783,  -18'd151,  
-18'd6157,  -18'd5094,  -18'd8168,  -18'd7285,  18'd202,  18'd4450,  -18'd3453,  18'd617,  -18'd1021,  -18'd1109,  -18'd102,  -18'd5766,  -18'd8516,  18'd5530,  -18'd6555,  18'd6453,  
-18'd7910,  18'd1009,  -18'd9801,  -18'd2782,  -18'd55,  18'd102,  -18'd1603,  -18'd903,  -18'd4133,  18'd5384,  -18'd558,  -18'd199,  -18'd4226,  -18'd2379,  18'd5749,  -18'd4089,  
-18'd2321,  18'd4652,  -18'd4758,  -18'd3674,  18'd7708,  18'd6765,  -18'd8423,  18'd3167,  -18'd6965,  -18'd7021,  -18'd9748,  18'd4418,  -18'd523,  -18'd2623,  18'd4639,  -18'd1712,  
18'd1295,  18'd8121,  18'd5285,  -18'd7589,  -18'd6124,  -18'd1854,  18'd4311,  18'd622,  18'd2561,  18'd1091,  -18'd7917,  -18'd4794,  -18'd7535,  18'd3129,  18'd2627,  18'd3517,  
18'd3141,  18'd1568,  -18'd3527,  -18'd3668,  -18'd7475,  -18'd6416,  18'd2110,  -18'd3017,  -18'd7729,  18'd4754,  18'd6615,  -18'd5798,  18'd1411,  -18'd5100,  -18'd4914,  -18'd3324,  
-18'd430,  18'd3635,  -18'd5502,  -18'd4468,  18'd6437,  -18'd4867,  -18'd7613,  -18'd6963,  18'd7148,  -18'd7780,  -18'd953,  -18'd4087,  18'd6410,  18'd3305,  18'd3348,  -18'd4963,  
-18'd6904,  -18'd724,  18'd2715,  -18'd1080,  -18'd6109,  -18'd3246,  -18'd3729,  18'd6051,  -18'd4339,  -18'd7709,  -18'd2505,  -18'd1089,  -18'd6925,  18'd4739,  -18'd894,  -18'd7848,  
18'd4429,  18'd5061,  -18'd78,  -18'd2264,  18'd456,  18'd2800,  18'd6976,  -18'd2357,  -18'd7494,  -18'd1101,  -18'd2040,  -18'd5550,  18'd8031,  -18'd6636,  -18'd3706,  18'd6233,  
-18'd6643,  -18'd6395,  -18'd7584,  18'd4641,  18'd6242,  -18'd531,  -18'd6232,  -18'd4982,  18'd8582,  -18'd7314,  18'd1639,  18'd5756,  18'd7188,  -18'd3650,  -18'd2752,  -18'd1811,  
18'd7058,  -18'd1112,  18'd6858,  -18'd7466,  18'd6131,  -18'd6503,  -18'd3476,  18'd714,  18'd7462,  -18'd9391,  -18'd2101,  -18'd8844,  -18'd74,  -18'd8358,  -18'd5416,  -18'd30,  
18'd4873,  -18'd9679,  18'd2134,  -18'd2774,  -18'd5238,  18'd4646,  -18'd163,  18'd318,  -18'd6563,  -18'd6500,  18'd5406,  18'd7495,  18'd2773,  -18'd8374,  -18'd6696,  18'd4964,  
-18'd8070,  -18'd5794,  18'd1040,  18'd1142,  -18'd1895,  18'd4388,  -18'd6749,  -18'd1656,  -18'd3984,  18'd3436,  -18'd932,  -18'd8421,  -18'd8882,  18'd4695,  -18'd7520,  -18'd6175,  

18'd9025,  18'd5534,  -18'd8869,  18'd787,  -18'd5883,  -18'd5174,  18'd8338,  18'd2078,  -18'd7568,  -18'd14099,  -18'd16558,  18'd706,  -18'd9061,  -18'd9094,  -18'd2685,  -18'd19589,  
18'd6565,  -18'd23440,  -18'd18228,  18'd14697,  -18'd2786,  -18'd4515,  -18'd2919,  -18'd5435,  -18'd15654,  18'd8288,  -18'd4287,  -18'd9886,  -18'd1668,  -18'd9626,  18'd14744,  -18'd21891,  
18'd10257,  18'd1332,  -18'd2066,  -18'd21617,  -18'd8111,  -18'd10434,  18'd20654,  18'd24826,  -18'd2152,  18'd13091,  -18'd12818,  18'd21079,  -18'd4702,  -18'd18911,  18'd17848,  -18'd14219,  
18'd16993,  18'd17315,  18'd9811,  -18'd24119,  -18'd5223,  18'd7201,  18'd1022,  18'd19108,  18'd14990,  -18'd17027,  18'd4829,  18'd10286,  -18'd4866,  -18'd1717,  18'd16782,  -18'd25801,  
18'd3483,  18'd15741,  18'd49,  18'd4301,  -18'd4175,  -18'd10952,  -18'd10612,  -18'd2161,  -18'd8187,  18'd1352,  -18'd6830,  -18'd1544,  -18'd8883,  18'd7842,  -18'd4146,  18'd6729,  
-18'd3568,  18'd1675,  -18'd5403,  18'd5604,  18'd6532,  -18'd15618,  -18'd13787,  18'd7173,  -18'd8541,  18'd20671,  -18'd2499,  18'd5560,  -18'd208,  18'd3358,  -18'd8434,  -18'd2001,  
18'd2152,  18'd17333,  -18'd7199,  -18'd5508,  -18'd5904,  18'd14482,  18'd5312,  18'd10949,  -18'd9718,  -18'd17821,  18'd9747,  18'd9181,  18'd3982,  18'd7008,  18'd11676,  18'd9877,  
-18'd2983,  18'd15890,  18'd15507,  -18'd1709,  18'd4042,  18'd305,  18'd2924,  18'd21027,  18'd1744,  18'd11539,  -18'd199,  18'd20828,  18'd6692,  -18'd3982,  18'd2862,  18'd26930,  
-18'd12269,  -18'd1114,  18'd4569,  -18'd28326,  18'd2281,  18'd2549,  -18'd8274,  -18'd4834,  -18'd3185,  -18'd5122,  -18'd13915,  18'd4261,  18'd5599,  18'd1885,  -18'd3396,  18'd15486,  
18'd896,  18'd7260,  -18'd6389,  18'd2275,  -18'd7703,  18'd9579,  -18'd2010,  -18'd18738,  18'd1753,  18'd7939,  -18'd1485,  18'd11094,  18'd2257,  18'd2347,  -18'd924,  -18'd13999,  
18'd9075,  -18'd84,  -18'd6031,  -18'd2696,  -18'd5306,  18'd2407,  -18'd13286,  18'd7198,  18'd7665,  18'd5301,  18'd14055,  18'd13078,  18'd4730,  18'd8137,  18'd1871,  -18'd4165,  
18'd6496,  -18'd933,  18'd29268,  18'd1426,  18'd4259,  -18'd10679,  18'd5772,  -18'd5007,  -18'd8418,  18'd20832,  18'd17612,  18'd6488,  18'd65,  18'd3346,  -18'd6294,  18'd7649,  
18'd6874,  -18'd11678,  18'd11475,  -18'd198,  -18'd1897,  18'd1476,  18'd14688,  18'd654,  -18'd214,  -18'd6384,  18'd20456,  -18'd4824,  -18'd4946,  18'd8868,  18'd11662,  18'd13423,  
18'd8060,  18'd11740,  18'd13446,  18'd7420,  -18'd3619,  18'd4918,  -18'd452,  -18'd20459,  18'd5147,  -18'd1403,  18'd5373,  -18'd12269,  18'd4284,  18'd13495,  -18'd4852,  18'd628,  
18'd11156,  18'd15851,  18'd2744,  18'd12136,  18'd5185,  -18'd4191,  -18'd2930,  -18'd4962,  18'd11039,  -18'd4835,  18'd3546,  -18'd10985,  -18'd3338,  -18'd734,  18'd4010,  18'd20445,  
-18'd976,  18'd8561,  -18'd10389,  18'd828,  18'd684,  -18'd2805,  18'd409,  -18'd4384,  18'd1874,  -18'd390,  -18'd194,  -18'd4682,  -18'd6916,  18'd2889,  18'd8282,  18'd2462,  

-18'd2280,  -18'd7974,  18'd5824,  -18'd6133,  -18'd4821,  18'd1657,  -18'd3547,  18'd5024,  18'd6958,  18'd1745,  18'd6652,  -18'd2116,  18'd7701,  -18'd7785,  -18'd4373,  18'd1949,  
18'd3383,  -18'd9396,  -18'd5818,  18'd1898,  18'd2408,  -18'd4042,  18'd7538,  -18'd8224,  -18'd1760,  -18'd7724,  -18'd7632,  18'd4790,  18'd6313,  18'd1884,  18'd4129,  -18'd7947,  
18'd1155,  18'd2992,  -18'd8376,  18'd7081,  -18'd1630,  18'd5183,  18'd4105,  -18'd1544,  -18'd2635,  18'd299,  -18'd9338,  -18'd506,  -18'd214,  18'd505,  -18'd3220,  -18'd1751,  
18'd5053,  18'd5343,  18'd146,  18'd5838,  -18'd2057,  -18'd9030,  -18'd1280,  18'd2776,  -18'd8686,  18'd4535,  -18'd1734,  -18'd7621,  18'd3476,  18'd1441,  -18'd7239,  18'd6715,  
-18'd9332,  18'd5973,  -18'd6150,  18'd8308,  18'd4172,  -18'd3143,  18'd6661,  -18'd580,  -18'd7586,  18'd5271,  18'd6484,  -18'd5794,  -18'd3708,  18'd1574,  -18'd5960,  -18'd5607,  
-18'd9019,  -18'd5217,  18'd6785,  -18'd2416,  18'd8270,  18'd4928,  18'd2738,  -18'd9869,  -18'd5447,  -18'd2756,  18'd5995,  -18'd7260,  18'd2217,  -18'd2863,  18'd5050,  18'd1798,  
-18'd5852,  18'd2829,  18'd5066,  -18'd4013,  -18'd5399,  -18'd2162,  -18'd628,  -18'd8510,  18'd3170,  -18'd8774,  18'd716,  18'd3256,  -18'd1490,  -18'd1923,  -18'd5662,  18'd4954,  
-18'd6729,  -18'd5591,  -18'd3488,  -18'd6372,  18'd364,  18'd7473,  -18'd8836,  18'd1949,  -18'd219,  -18'd5243,  18'd2177,  -18'd4780,  18'd5429,  18'd3265,  -18'd3983,  -18'd8582,  
-18'd4259,  18'd1411,  18'd5019,  -18'd4397,  18'd3233,  18'd5479,  -18'd5675,  -18'd1755,  18'd140,  -18'd945,  -18'd1261,  -18'd967,  -18'd8645,  -18'd8776,  18'd6025,  -18'd1816,  
-18'd5287,  18'd5982,  18'd5569,  18'd2471,  -18'd7655,  -18'd1427,  -18'd2514,  18'd5861,  18'd3409,  -18'd6454,  -18'd6932,  -18'd8220,  18'd565,  18'd5389,  -18'd8182,  -18'd3296,  
-18'd2345,  -18'd10691,  18'd3236,  -18'd9767,  -18'd4202,  -18'd2010,  -18'd9201,  -18'd6869,  -18'd9532,  18'd2156,  -18'd3422,  -18'd10693,  18'd746,  -18'd3270,  -18'd4298,  -18'd7205,  
18'd2081,  -18'd10266,  18'd4841,  18'd6934,  18'd7406,  18'd5604,  -18'd7537,  18'd483,  -18'd3556,  -18'd5283,  18'd5168,  -18'd7122,  -18'd7549,  18'd3066,  -18'd8169,  18'd2288,  
18'd210,  -18'd1774,  18'd1806,  18'd3256,  18'd1622,  -18'd7577,  18'd4614,  -18'd3689,  18'd5943,  18'd3562,  18'd6399,  18'd3565,  -18'd5106,  18'd766,  18'd6243,  18'd5984,  
-18'd7830,  -18'd11263,  -18'd172,  -18'd4795,  18'd6053,  -18'd8865,  -18'd4952,  18'd474,  18'd6156,  18'd3769,  18'd871,  -18'd9534,  18'd7879,  -18'd9141,  18'd6718,  -18'd4171,  
-18'd6451,  -18'd9214,  -18'd2718,  -18'd5809,  -18'd1383,  -18'd8441,  18'd850,  18'd4693,  -18'd9338,  18'd6113,  18'd2531,  -18'd4303,  -18'd3517,  18'd1364,  18'd5240,  -18'd10599,  
18'd4367,  -18'd8342,  -18'd6507,  18'd5445,  -18'd520,  18'd2701,  -18'd8739,  -18'd8130,  -18'd687,  -18'd2140,  18'd1720,  -18'd5364,  18'd3920,  -18'd8422,  -18'd5467,  18'd872,  

-18'd1336,  18'd3238,  -18'd12256,  18'd1844,  -18'd2832,  -18'd8300,  -18'd4082,  -18'd141,  -18'd59,  -18'd12599,  18'd4817,  18'd4234,  18'd8556,  -18'd2379,  -18'd11758,  -18'd2113,  
-18'd9416,  -18'd10495,  -18'd847,  18'd3432,  18'd25,  -18'd4699,  18'd1452,  -18'd3007,  18'd4882,  -18'd3402,  -18'd1811,  -18'd5308,  18'd4377,  18'd1535,  -18'd9249,  -18'd11490,  
-18'd3158,  -18'd5078,  18'd599,  -18'd4802,  18'd3045,  -18'd1553,  -18'd4653,  18'd2148,  18'd1385,  -18'd2207,  -18'd7846,  -18'd8454,  -18'd1136,  18'd2019,  18'd461,  18'd3386,  
18'd413,  -18'd2331,  18'd2148,  -18'd396,  -18'd1962,  -18'd318,  -18'd4189,  -18'd3570,  -18'd3629,  18'd4038,  -18'd9645,  18'd2492,  18'd4020,  -18'd9379,  -18'd2435,  18'd2491,  
-18'd7680,  18'd5772,  18'd1150,  18'd4511,  18'd7141,  -18'd8114,  18'd1918,  -18'd1438,  -18'd9756,  -18'd3871,  18'd1659,  -18'd8702,  18'd8744,  -18'd4890,  18'd2331,  18'd8551,  
-18'd1480,  -18'd7356,  18'd920,  18'd648,  18'd6626,  -18'd241,  -18'd11574,  -18'd9585,  18'd1594,  18'd2688,  18'd4717,  -18'd7879,  -18'd904,  -18'd1846,  -18'd4899,  -18'd3412,  
18'd4715,  18'd2419,  18'd87,  -18'd3180,  18'd7008,  -18'd1496,  18'd1557,  18'd888,  -18'd4384,  -18'd10996,  -18'd9360,  -18'd2738,  18'd4282,  18'd499,  18'd6768,  -18'd192,  
18'd1715,  -18'd6426,  18'd383,  -18'd9433,  -18'd1706,  -18'd6064,  18'd2638,  -18'd2421,  -18'd742,  -18'd9318,  -18'd749,  -18'd9271,  18'd8915,  -18'd10664,  -18'd8513,  -18'd581,  
18'd272,  -18'd7664,  -18'd4722,  -18'd8760,  -18'd8791,  -18'd9346,  -18'd7113,  -18'd6547,  18'd6580,  -18'd1021,  18'd2718,  -18'd424,  -18'd20,  -18'd6937,  -18'd12209,  -18'd7166,  
-18'd884,  18'd7295,  18'd2441,  -18'd899,  18'd4085,  18'd4302,  18'd2582,  -18'd6709,  18'd3516,  -18'd829,  18'd2695,  -18'd2788,  18'd7526,  18'd4757,  -18'd9850,  -18'd2840,  
18'd3598,  -18'd10389,  -18'd9009,  -18'd2217,  18'd5249,  18'd2865,  -18'd3943,  18'd7647,  -18'd3072,  -18'd2785,  -18'd9258,  18'd734,  -18'd816,  18'd4861,  -18'd11575,  18'd2021,  
-18'd4138,  -18'd2187,  -18'd7979,  -18'd12361,  18'd1344,  18'd2152,  -18'd7292,  -18'd9619,  -18'd1700,  -18'd1190,  -18'd9633,  -18'd172,  18'd2410,  -18'd9872,  -18'd8797,  -18'd6598,  
-18'd4882,  -18'd6664,  -18'd9604,  -18'd3840,  18'd5410,  -18'd6316,  -18'd862,  18'd2066,  18'd2583,  -18'd4485,  -18'd891,  -18'd5551,  -18'd1423,  -18'd9476,  18'd1239,  18'd7096,  
-18'd6230,  18'd3520,  -18'd7008,  -18'd7630,  -18'd8264,  -18'd5257,  -18'd6875,  18'd1788,  18'd1177,  18'd2773,  18'd869,  -18'd7797,  -18'd7264,  18'd2487,  -18'd9693,  18'd655,  
-18'd3352,  18'd6628,  -18'd3429,  -18'd2472,  -18'd2475,  18'd3359,  -18'd720,  -18'd5152,  18'd2638,  -18'd4626,  -18'd3614,  18'd5337,  18'd737,  18'd1235,  18'd2530,  -18'd4199,  
-18'd1067,  18'd724,  -18'd8331,  -18'd5927,  18'd1669,  -18'd5144,  -18'd9091,  18'd8169,  -18'd827,  -18'd1757,  18'd3889,  18'd2846,  -18'd4469,  -18'd11063,  -18'd155,  -18'd6553,  

18'd15620,  -18'd5035,  18'd11042,  18'd20961,  18'd1846,  18'd4598,  18'd1340,  -18'd1887,  -18'd2149,  18'd6081,  -18'd2819,  18'd6420,  -18'd2978,  18'd2084,  -18'd17750,  18'd16364,  
-18'd9287,  18'd5205,  18'd7075,  -18'd3777,  18'd6137,  -18'd5562,  18'd2775,  -18'd8945,  -18'd3082,  -18'd7532,  18'd3211,  -18'd5628,  18'd7982,  18'd12931,  -18'd11105,  18'd5187,  
-18'd6735,  18'd13386,  18'd11457,  -18'd8079,  -18'd7812,  -18'd8089,  18'd896,  -18'd8618,  18'd4155,  -18'd5514,  -18'd5550,  18'd8576,  -18'd2060,  18'd7633,  -18'd13652,  18'd14192,  
-18'd18288,  18'd11629,  -18'd5243,  -18'd2714,  -18'd3852,  18'd5076,  18'd12072,  -18'd4787,  -18'd6166,  18'd867,  -18'd3631,  18'd10969,  -18'd1166,  18'd18037,  -18'd20998,  18'd8457,  
18'd11003,  -18'd10379,  18'd9366,  18'd24768,  -18'd2272,  18'd12174,  -18'd5287,  18'd814,  18'd3770,  18'd21462,  18'd190,  18'd21359,  -18'd5276,  18'd4068,  -18'd1646,  -18'd1553,  
-18'd2497,  -18'd4588,  -18'd2232,  18'd5136,  18'd6189,  -18'd7060,  -18'd17664,  18'd2470,  18'd11689,  18'd6465,  18'd18897,  18'd7265,  18'd6683,  18'd9510,  -18'd2460,  -18'd5331,  
18'd2043,  -18'd520,  -18'd19363,  -18'd1356,  18'd5868,  -18'd6220,  -18'd32065,  -18'd10725,  -18'd4909,  18'd13391,  18'd18032,  18'd25034,  18'd5048,  -18'd917,  18'd11828,  18'd7390,  
18'd2497,  18'd4678,  -18'd14911,  -18'd14043,  -18'd8957,  -18'd11673,  -18'd8399,  18'd2295,  18'd9300,  18'd23523,  -18'd12383,  18'd13833,  18'd6720,  18'd3367,  18'd9490,  18'd10223,  
18'd1796,  -18'd6958,  18'd3440,  -18'd10167,  18'd5715,  -18'd5125,  -18'd4218,  -18'd12039,  -18'd245,  18'd4751,  -18'd2226,  18'd8180,  18'd6184,  18'd11196,  -18'd3172,  18'd3266,  
-18'd8704,  -18'd7635,  18'd11967,  -18'd8807,  18'd3191,  -18'd7292,  18'd4666,  -18'd5878,  -18'd1887,  18'd12604,  18'd1397,  18'd14510,  18'd1267,  18'd3536,  -18'd4273,  -18'd4201,  
-18'd2283,  -18'd6019,  -18'd23047,  -18'd1038,  -18'd14,  -18'd6878,  18'd1720,  18'd1180,  18'd4859,  18'd4005,  18'd2991,  -18'd5663,  -18'd1530,  -18'd3296,  18'd3120,  -18'd1909,  
-18'd2341,  -18'd13006,  -18'd10073,  18'd2622,  -18'd4109,  -18'd23688,  -18'd2658,  18'd3537,  -18'd1751,  18'd16305,  18'd12157,  18'd1500,  18'd928,  -18'd17255,  18'd10933,  18'd14240,  
-18'd569,  -18'd7282,  -18'd5333,  -18'd9729,  -18'd7734,  18'd265,  18'd12395,  18'd11368,  -18'd6462,  18'd1977,  18'd20916,  18'd4117,  18'd3297,  -18'd11404,  18'd798,  18'd6977,  
-18'd7592,  -18'd14294,  18'd3983,  -18'd280,  -18'd2074,  18'd4261,  18'd17028,  18'd9043,  18'd535,  18'd6565,  18'd7622,  -18'd2691,  18'd2063,  -18'd2969,  18'd4392,  18'd561,  
18'd4798,  -18'd19530,  -18'd7544,  18'd6027,  18'd5358,  18'd2949,  18'd19194,  -18'd28095,  18'd405,  -18'd1733,  18'd6975,  -18'd53,  18'd5802,  -18'd15117,  18'd16820,  -18'd17443,  
18'd9658,  -18'd35707,  18'd9238,  -18'd2930,  -18'd7005,  -18'd29042,  18'd8752,  -18'd179,  -18'd490,  -18'd1237,  -18'd17390,  -18'd19298,  18'd2110,  -18'd26700,  18'd19676,  -18'd4464,  

-18'd16503,  18'd19357,  18'd4547,  18'd11711,  -18'd3456,  -18'd1317,  18'd15119,  18'd992,  18'd5034,  -18'd2863,  18'd14277,  -18'd5048,  -18'd1457,  18'd4765,  -18'd10155,  18'd6763,  
18'd470,  18'd6008,  18'd8467,  -18'd1758,  -18'd4338,  18'd6479,  -18'd5173,  18'd4195,  -18'd9251,  18'd9668,  18'd9540,  18'd13208,  18'd4751,  18'd4495,  -18'd7705,  18'd7477,  
-18'd11438,  18'd21091,  18'd9117,  -18'd3129,  18'd8071,  18'd11854,  -18'd14150,  18'd11612,  18'd11071,  18'd7103,  18'd798,  18'd15012,  -18'd3542,  18'd16432,  -18'd22716,  18'd20287,  
-18'd6357,  18'd11562,  -18'd2228,  18'd25727,  -18'd3897,  -18'd13547,  -18'd21225,  -18'd17555,  -18'd6413,  -18'd1061,  -18'd19014,  -18'd997,  18'd9447,  18'd4520,  -18'd12983,  18'd25991,  
-18'd161,  -18'd767,  -18'd144,  18'd2176,  -18'd7113,  -18'd3947,  18'd1607,  18'd1037,  18'd1153,  18'd1829,  -18'd6928,  -18'd7627,  18'd4325,  18'd5739,  18'd3050,  18'd5978,  
18'd7823,  -18'd4050,  -18'd11577,  -18'd6568,  18'd2887,  18'd5933,  -18'd16413,  -18'd10421,  -18'd2631,  -18'd5139,  -18'd2910,  18'd3814,  18'd1362,  -18'd359,  -18'd6092,  18'd7765,  
18'd3417,  -18'd3467,  -18'd10955,  -18'd3464,  18'd504,  18'd12414,  -18'd13742,  -18'd15801,  -18'd1184,  18'd10234,  -18'd149,  -18'd1435,  18'd7433,  18'd17714,  18'd12818,  18'd11073,  
-18'd4468,  -18'd6606,  -18'd16390,  18'd7913,  -18'd6800,  -18'd10975,  -18'd16738,  -18'd10473,  -18'd6119,  18'd18032,  -18'd9194,  18'd682,  18'd6686,  -18'd93,  18'd17688,  18'd181,  
18'd14084,  -18'd23057,  -18'd2493,  -18'd1248,  -18'd7729,  -18'd8381,  18'd1436,  -18'd8347,  18'd5313,  18'd9403,  -18'd11993,  18'd2458,  18'd8185,  18'd11865,  18'd8139,  -18'd10653,  
18'd581,  -18'd6670,  -18'd13358,  18'd5503,  -18'd6403,  -18'd15214,  -18'd2854,  -18'd5881,  -18'd8245,  18'd2678,  -18'd1633,  -18'd9408,  -18'd716,  -18'd6056,  18'd15955,  -18'd5072,  
-18'd2538,  -18'd408,  18'd9871,  -18'd5227,  -18'd570,  -18'd6530,  18'd3400,  18'd72,  18'd2007,  -18'd3608,  18'd5711,  -18'd5875,  18'd731,  -18'd8925,  18'd1254,  -18'd8166,  
18'd641,  18'd10233,  -18'd7251,  -18'd4263,  18'd7075,  18'd11889,  18'd6228,  18'd7978,  -18'd4264,  18'd6056,  -18'd6394,  -18'd3641,  18'd9047,  18'd9890,  18'd5327,  18'd9882,  
18'd8581,  -18'd10655,  -18'd22783,  18'd12860,  18'd4420,  -18'd3966,  -18'd461,  18'd16975,  -18'd15016,  18'd9791,  18'd10080,  18'd704,  -18'd3676,  -18'd910,  18'd15790,  -18'd14719,  
-18'd12592,  -18'd9472,  18'd9612,  18'd4687,  18'd3682,  -18'd4907,  -18'd750,  18'd13795,  -18'd9154,  18'd4871,  18'd4320,  -18'd8992,  -18'd3527,  18'd516,  18'd8326,  -18'd12481,  
18'd3621,  -18'd2142,  18'd7728,  -18'd13256,  -18'd3557,  -18'd6093,  18'd8043,  18'd1247,  -18'd10802,  18'd10782,  18'd4321,  18'd3587,  18'd4521,  -18'd11181,  18'd14244,  -18'd6786,  
-18'd2406,  -18'd764,  18'd16369,  18'd6429,  18'd2870,  18'd4805,  18'd8280,  18'd4891,  -18'd4818,  -18'd10313,  18'd7228,  18'd4811,  -18'd1202,  -18'd8229,  18'd3880,  18'd1082,  

-18'd27928,  18'd13105,  18'd23622,  -18'd11411,  -18'd3208,  18'd8043,  18'd10682,  18'd2690,  18'd3190,  -18'd13699,  -18'd2300,  -18'd28141,  -18'd1451,  -18'd11040,  -18'd2691,  18'd22146,  
-18'd13035,  -18'd3688,  -18'd3314,  18'd13856,  18'd2617,  18'd2796,  18'd11487,  18'd8103,  -18'd1363,  -18'd5223,  -18'd4949,  18'd886,  -18'd2980,  18'd5914,  18'd3407,  18'd4874,  
18'd6431,  18'd9518,  -18'd2159,  18'd16629,  -18'd1868,  18'd11661,  18'd4184,  18'd1192,  -18'd16053,  -18'd18093,  -18'd18224,  -18'd16248,  18'd3364,  18'd11963,  -18'd8590,  -18'd3017,  
-18'd10000,  18'd28159,  -18'd9595,  -18'd4266,  18'd4846,  18'd9252,  -18'd10616,  18'd4951,  -18'd7280,  -18'd4981,  -18'd22456,  18'd9297,  18'd3407,  18'd19631,  -18'd11766,  18'd5008,  
-18'd8003,  18'd4246,  18'd8859,  18'd705,  18'd7719,  -18'd5283,  -18'd5908,  18'd12996,  -18'd4526,  -18'd2352,  18'd1464,  -18'd10977,  18'd11039,  18'd3443,  18'd662,  18'd18736,  
-18'd9002,  -18'd16311,  18'd1234,  18'd13221,  -18'd4205,  18'd8561,  18'd12737,  -18'd13528,  -18'd9169,  18'd5055,  18'd10384,  18'd2152,  18'd222,  18'd7710,  18'd10266,  18'd5983,  
18'd190,  18'd2519,  -18'd11388,  18'd4252,  18'd8263,  18'd15830,  -18'd17851,  -18'd2255,  -18'd10877,  18'd6911,  -18'd2381,  18'd1272,  18'd3760,  18'd8290,  -18'd12376,  18'd22,  
-18'd7447,  -18'd839,  -18'd17732,  -18'd3150,  18'd3924,  -18'd3977,  -18'd11345,  18'd1934,  18'd10544,  18'd2581,  -18'd11034,  -18'd954,  -18'd456,  18'd8979,  18'd13616,  18'd10601,  
-18'd14490,  -18'd10816,  -18'd6537,  -18'd755,  18'd2205,  -18'd6994,  -18'd4607,  18'd10268,  -18'd7127,  18'd14015,  -18'd16749,  -18'd4089,  -18'd4113,  -18'd3581,  -18'd754,  -18'd5505,  
-18'd6015,  -18'd13996,  18'd7966,  -18'd16424,  -18'd526,  -18'd3069,  -18'd9701,  18'd19054,  -18'd10737,  18'd19513,  18'd8813,  18'd14343,  18'd5414,  18'd10322,  18'd595,  -18'd1007,  
18'd888,  -18'd6383,  18'd79,  18'd5763,  -18'd934,  -18'd3984,  -18'd20056,  18'd14974,  -18'd5613,  18'd9776,  -18'd3209,  18'd18041,  -18'd2414,  18'd1229,  18'd6663,  18'd12559,  
18'd11823,  -18'd16684,  -18'd17203,  18'd8742,  -18'd542,  18'd2038,  18'd12080,  -18'd10314,  18'd8402,  -18'd12033,  18'd852,  18'd10561,  -18'd306,  18'd1319,  18'd6679,  18'd4824,  
-18'd36538,  18'd1322,  -18'd2530,  18'd5054,  18'd2690,  -18'd2467,  -18'd4779,  18'd4772,  -18'd23457,  18'd26151,  -18'd9925,  -18'd7667,  18'd6781,  18'd2160,  18'd4455,  -18'd2498,  
-18'd20753,  -18'd9399,  18'd10506,  -18'd3395,  18'd2955,  -18'd4619,  18'd1,  18'd34905,  -18'd12094,  18'd29437,  18'd17083,  -18'd6283,  -18'd1242,  -18'd4988,  18'd12085,  18'd6256,  
-18'd8310,  -18'd7323,  18'd5550,  18'd13066,  -18'd8102,  -18'd11618,  -18'd1850,  18'd649,  -18'd957,  18'd1717,  18'd11633,  18'd9096,  18'd5113,  18'd7376,  18'd11905,  -18'd8796,  
18'd8843,  -18'd9563,  18'd2004,  18'd3220,  18'd4971,  -18'd12236,  18'd3205,  18'd4962,  18'd15415,  -18'd13747,  -18'd4158,  -18'd2387,  18'd3749,  -18'd12308,  18'd18551,  -18'd9292,  

-18'd18699,  18'd379,  18'd12461,  18'd9438,  -18'd5970,  -18'd11305,  18'd6025,  18'd6511,  -18'd10367,  -18'd15770,  -18'd8854,  -18'd14123,  18'd1379,  -18'd4610,  -18'd10955,  -18'd17549,  
-18'd17292,  18'd943,  18'd7741,  -18'd17652,  -18'd3809,  -18'd18373,  18'd1062,  -18'd11137,  -18'd6286,  -18'd4418,  -18'd6914,  -18'd11805,  18'd715,  -18'd3537,  -18'd6593,  -18'd12539,  
-18'd7270,  -18'd3815,  -18'd9064,  -18'd14883,  -18'd3903,  -18'd752,  -18'd411,  -18'd10495,  -18'd6930,  -18'd7519,  -18'd8040,  18'd5959,  18'd1712,  -18'd9377,  -18'd2477,  -18'd10183,  
18'd20379,  -18'd1453,  -18'd5744,  -18'd22077,  18'd3396,  18'd28772,  18'd1443,  -18'd10356,  18'd24089,  18'd1307,  -18'd15497,  -18'd16014,  -18'd4734,  18'd11653,  18'd11480,  -18'd14112,  
-18'd21074,  18'd7634,  18'd1766,  18'd20209,  -18'd3305,  -18'd15058,  18'd3480,  18'd16348,  -18'd7683,  18'd16162,  18'd435,  18'd2899,  18'd3019,  18'd17705,  18'd1077,  18'd5150,  
-18'd10106,  18'd19401,  -18'd15127,  18'd9965,  -18'd7624,  -18'd3919,  -18'd997,  18'd8568,  18'd2050,  -18'd3567,  -18'd14185,  -18'd21260,  18'd2520,  -18'd2518,  -18'd16147,  18'd12840,  
-18'd3643,  18'd244,  18'd1803,  18'd18952,  -18'd6870,  -18'd7082,  18'd2577,  18'd10914,  -18'd4170,  -18'd6702,  18'd4140,  -18'd4130,  18'd9403,  18'd9750,  -18'd14136,  18'd8547,  
18'd4446,  -18'd19812,  18'd3141,  18'd1078,  18'd2917,  18'd12387,  18'd10121,  18'd2701,  18'd15787,  -18'd5328,  -18'd1947,  -18'd6022,  -18'd2921,  18'd3054,  18'd6031,  18'd2658,  
-18'd20971,  18'd4110,  -18'd7748,  18'd12699,  18'd777,  -18'd10231,  -18'd5922,  18'd17959,  -18'd706,  18'd18961,  -18'd17128,  18'd16572,  18'd10235,  18'd4276,  -18'd7669,  18'd2456,  
-18'd2399,  18'd2782,  -18'd18718,  18'd8955,  18'd4177,  18'd5546,  18'd1686,  -18'd12945,  -18'd10857,  18'd1795,  18'd15394,  18'd18878,  18'd3175,  18'd1825,  -18'd2203,  -18'd3723,  
-18'd1645,  18'd22942,  18'd8514,  18'd13932,  18'd7478,  -18'd4830,  18'd6375,  18'd2039,  -18'd730,  18'd3098,  -18'd545,  18'd3345,  18'd8396,  18'd9430,  18'd13296,  18'd6091,  
18'd3587,  18'd2132,  18'd17054,  -18'd3276,  -18'd731,  -18'd3535,  18'd5433,  18'd361,  18'd4117,  18'd4269,  18'd2352,  18'd3443,  -18'd1071,  18'd2634,  18'd6991,  18'd4030,  
18'd3659,  -18'd26664,  -18'd11987,  18'd6725,  -18'd3705,  -18'd2372,  18'd4526,  -18'd15567,  -18'd6128,  18'd5906,  18'd7221,  -18'd2652,  18'd6672,  -18'd5198,  18'd19956,  -18'd16812,  
18'd2047,  -18'd1332,  -18'd7099,  18'd1270,  18'd3319,  -18'd1585,  -18'd2624,  -18'd7053,  -18'd4585,  -18'd5915,  18'd13432,  18'd3351,  -18'd3696,  -18'd5414,  18'd15444,  18'd2771,  
18'd10321,  18'd2177,  18'd3088,  -18'd2358,  -18'd3166,  18'd597,  18'd2053,  -18'd10595,  18'd10333,  -18'd247,  18'd11054,  18'd12286,  18'd9575,  18'd4709,  18'd21184,  -18'd6929,  
-18'd4230,  18'd28339,  18'd10504,  -18'd13680,  18'd107,  -18'd1583,  -18'd6102,  -18'd745,  18'd17387,  18'd8224,  18'd9107,  18'd2082,  -18'd2776,  18'd1025,  18'd7508,  18'd16807,  

18'd1478,  -18'd4224,  -18'd3362,  -18'd392,  18'd6616,  18'd6047,  18'd2120,  18'd7259,  18'd4469,  -18'd7699,  -18'd9512,  18'd447,  18'd106,  18'd6565,  18'd6361,  -18'd7221,  
18'd6942,  -18'd9684,  -18'd6120,  -18'd6002,  18'd1411,  -18'd2452,  -18'd198,  -18'd6461,  -18'd5305,  18'd1465,  -18'd8786,  18'd1598,  -18'd5750,  18'd3301,  -18'd8882,  -18'd2623,  
-18'd3514,  18'd764,  18'd1611,  18'd254,  18'd1765,  -18'd1677,  18'd559,  18'd5594,  -18'd11075,  -18'd9905,  18'd5762,  -18'd2200,  -18'd516,  -18'd6249,  -18'd7234,  -18'd6249,  
-18'd4754,  18'd895,  -18'd5841,  -18'd10471,  -18'd71,  18'd4331,  -18'd3944,  18'd6469,  18'd4688,  -18'd8632,  -18'd7754,  -18'd6777,  18'd7776,  -18'd8881,  -18'd11234,  18'd1273,  
18'd1788,  18'd2614,  18'd2116,  18'd1830,  -18'd2540,  18'd976,  18'd254,  -18'd7076,  -18'd3776,  -18'd5831,  18'd2298,  -18'd10173,  -18'd5828,  18'd1751,  -18'd2616,  18'd3538,  
18'd776,  -18'd6427,  18'd659,  18'd7701,  18'd7410,  18'd2834,  -18'd3884,  18'd7779,  -18'd461,  18'd373,  -18'd7932,  -18'd4640,  18'd7929,  -18'd4917,  -18'd3548,  -18'd6026,  
18'd4240,  -18'd7308,  -18'd4954,  -18'd3582,  18'd296,  -18'd3958,  -18'd3948,  -18'd8450,  18'd4045,  -18'd8974,  18'd2799,  -18'd6160,  -18'd7596,  -18'd10000,  -18'd2027,  18'd2226,  
18'd4984,  -18'd4965,  -18'd8570,  18'd5779,  -18'd6136,  -18'd4700,  18'd3665,  -18'd2554,  -18'd7605,  18'd1284,  18'd160,  -18'd9513,  -18'd6144,  -18'd6686,  -18'd8286,  -18'd1543,  
-18'd4960,  -18'd8870,  -18'd3168,  18'd2189,  -18'd4286,  -18'd7674,  -18'd7247,  18'd3550,  18'd831,  -18'd1042,  18'd4091,  18'd3820,  18'd1881,  18'd6907,  -18'd6598,  -18'd4131,  
-18'd8208,  -18'd4854,  -18'd3575,  -18'd5989,  18'd1641,  -18'd156,  18'd4022,  -18'd7100,  -18'd2043,  18'd492,  18'd5412,  -18'd240,  -18'd7444,  18'd2003,  -18'd1540,  -18'd5628,  
-18'd820,  18'd4630,  18'd3478,  18'd2037,  -18'd1501,  -18'd4707,  18'd975,  18'd6600,  -18'd8368,  -18'd9080,  18'd5029,  -18'd2110,  18'd3915,  18'd6863,  18'd1247,  18'd897,  
18'd3263,  18'd394,  18'd2771,  18'd1190,  18'd2130,  -18'd4471,  18'd4750,  18'd2660,  18'd1281,  18'd3686,  -18'd1810,  -18'd7960,  -18'd3143,  -18'd3451,  18'd209,  18'd1432,  
18'd5631,  -18'd2827,  -18'd2510,  18'd3669,  -18'd5925,  -18'd10656,  -18'd4084,  -18'd5716,  18'd4980,  -18'd4952,  18'd1929,  -18'd7051,  18'd7068,  -18'd5677,  -18'd4130,  -18'd2208,  
18'd690,  18'd1075,  -18'd7593,  18'd672,  18'd5697,  -18'd10586,  -18'd8787,  -18'd1514,  -18'd9343,  -18'd1365,  18'd2412,  18'd3294,  18'd244,  -18'd416,  -18'd11030,  -18'd7827,  
18'd3821,  18'd5060,  -18'd9799,  -18'd2141,  18'd464,  18'd4066,  18'd1462,  -18'd6228,  18'd1334,  18'd4676,  18'd2750,  -18'd2492,  -18'd5152,  18'd6188,  -18'd6593,  -18'd8100,  
-18'd5132,  18'd3783,  18'd6047,  18'd4690,  -18'd4804,  -18'd1439,  18'd3011,  -18'd8326,  -18'd9059,  -18'd2794,  -18'd4316,  -18'd9542,  -18'd1320,  -18'd8029,  -18'd2559,  18'd2590,  

18'd11814,  18'd16515,  18'd6877,  18'd22534,  -18'd6438,  18'd8815,  -18'd2636,  18'd3955,  18'd1039,  -18'd12221,  -18'd7442,  -18'd9603,  -18'd1559,  -18'd1291,  -18'd3683,  18'd17490,  
-18'd16182,  18'd19973,  18'd13643,  -18'd9735,  18'd8267,  18'd1107,  -18'd1438,  18'd3275,  18'd4860,  -18'd18166,  18'd2317,  -18'd20738,  -18'd1962,  18'd5702,  -18'd7649,  18'd9953,  
-18'd14456,  18'd21508,  -18'd537,  18'd8256,  18'd3397,  -18'd979,  -18'd3320,  18'd13211,  -18'd8374,  -18'd5830,  -18'd13483,  -18'd28998,  -18'd6567,  -18'd20433,  18'd4891,  18'd14630,  
18'd6928,  -18'd12295,  -18'd30433,  18'd765,  -18'd3823,  -18'd26660,  18'd16843,  18'd4488,  -18'd12108,  -18'd9955,  -18'd24607,  -18'd40383,  -18'd4615,  -18'd13409,  18'd6225,  -18'd12725,  
18'd5220,  -18'd3186,  -18'd7199,  18'd7870,  18'd8423,  18'd13290,  18'd145,  18'd5082,  18'd11304,  18'd2644,  18'd8868,  -18'd3558,  18'd6357,  18'd6287,  18'd2633,  -18'd4089,  
-18'd11595,  -18'd4404,  18'd11115,  18'd2645,  18'd1158,  -18'd2445,  -18'd1637,  -18'd115,  18'd13545,  -18'd15726,  -18'd3507,  18'd1224,  -18'd10234,  18'd779,  18'd6752,  18'd3895,  
-18'd3950,  18'd3579,  -18'd2053,  18'd18629,  18'd4393,  -18'd15976,  18'd9524,  -18'd8756,  18'd7562,  18'd10438,  -18'd14406,  -18'd17102,  18'd2631,  -18'd320,  18'd6442,  18'd15746,  
-18'd1678,  -18'd23263,  -18'd15460,  18'd2399,  18'd880,  -18'd13653,  -18'd7931,  -18'd8047,  -18'd15943,  -18'd2435,  -18'd13374,  -18'd8326,  -18'd10374,  -18'd6674,  18'd1769,  -18'd14134,  
18'd4867,  -18'd13788,  18'd2793,  18'd6121,  18'd4596,  18'd8290,  18'd15129,  18'd3471,  -18'd5468,  18'd9443,  18'd11418,  -18'd3275,  -18'd8194,  -18'd1394,  18'd6381,  -18'd12122,  
-18'd854,  18'd3827,  18'd8207,  18'd8734,  18'd121,  18'd14337,  18'd17508,  18'd9122,  18'd17230,  -18'd10671,  18'd4366,  -18'd11995,  -18'd1447,  -18'd8129,  -18'd6593,  -18'd9252,  
18'd9731,  -18'd10513,  18'd6605,  18'd1030,  18'd4325,  18'd10411,  18'd9577,  -18'd19474,  -18'd6871,  -18'd3297,  18'd7096,  -18'd3413,  -18'd708,  18'd7784,  -18'd10624,  18'd13885,  
18'd5753,  -18'd16046,  -18'd1814,  18'd5437,  -18'd1541,  -18'd7672,  -18'd10671,  -18'd15502,  -18'd19181,  18'd5150,  -18'd8554,  -18'd9162,  -18'd6804,  18'd706,  -18'd8821,  -18'd11811,  
18'd12280,  18'd15344,  18'd7178,  -18'd1304,  -18'd4518,  18'd623,  18'd2658,  -18'd3728,  18'd6465,  18'd635,  18'd8254,  18'd9005,  18'd2776,  18'd4903,  -18'd6814,  -18'd18176,  
-18'd12552,  18'd2664,  18'd4139,  18'd11409,  18'd5864,  18'd15470,  -18'd9968,  18'd6837,  18'd16239,  -18'd15644,  -18'd11503,  18'd13562,  -18'd5058,  18'd1151,  18'd553,  18'd7193,  
18'd14396,  -18'd597,  18'd7750,  -18'd11486,  18'd5959,  18'd15801,  18'd13301,  18'd1666,  -18'd5513,  18'd8079,  -18'd1000,  18'd25859,  18'd1074,  18'd936,  -18'd7347,  18'd5112,  
18'd7647,  18'd8039,  18'd21463,  18'd1430,  18'd2865,  18'd8153,  -18'd8575,  -18'd7522,  18'd3856,  18'd10576,  18'd4680,  18'd3457,  -18'd4075,  18'd23809,  18'd69,  18'd9827,  

18'd3140,  -18'd1198,  -18'd9277,  18'd6379,  -18'd4496,  -18'd6537,  -18'd13036,  18'd1578,  18'd4319,  18'd13487,  -18'd14813,  18'd4293,  -18'd4804,  18'd3934,  -18'd356,  18'd6576,  
-18'd6497,  -18'd11857,  -18'd5921,  18'd8491,  -18'd6669,  -18'd8732,  -18'd8706,  -18'd10243,  18'd3657,  -18'd5720,  -18'd5992,  18'd2986,  18'd6640,  -18'd925,  -18'd7999,  18'd735,  
-18'd7190,  18'd4640,  -18'd6518,  -18'd5336,  -18'd8304,  -18'd4295,  -18'd407,  -18'd8114,  -18'd5216,  18'd752,  -18'd58,  -18'd2906,  -18'd1234,  -18'd2567,  -18'd4905,  18'd2741,  
-18'd5007,  18'd4973,  18'd6233,  18'd3661,  18'd8535,  18'd4193,  -18'd3762,  -18'd6235,  -18'd12080,  18'd4698,  -18'd949,  -18'd7144,  18'd7154,  18'd2898,  -18'd12235,  -18'd12704,  
-18'd9042,  18'd928,  18'd2824,  -18'd3377,  18'd2397,  18'd430,  18'd2460,  18'd654,  -18'd10419,  18'd7021,  -18'd13427,  -18'd3820,  18'd3346,  18'd476,  -18'd6010,  -18'd2930,  
18'd7316,  -18'd13128,  18'd3223,  -18'd6068,  -18'd2747,  -18'd11806,  -18'd4306,  18'd159,  -18'd6214,  18'd9598,  -18'd4349,  -18'd1945,  18'd141,  -18'd3980,  -18'd2225,  -18'd10998,  
-18'd194,  -18'd8065,  18'd4745,  -18'd5335,  18'd8697,  18'd1412,  -18'd8166,  -18'd1417,  -18'd1798,  18'd7375,  18'd751,  -18'd10510,  -18'd5959,  -18'd2691,  -18'd8830,  -18'd449,  
18'd925,  18'd4886,  -18'd5503,  18'd2881,  -18'd6296,  -18'd4802,  18'd5427,  -18'd10027,  -18'd9135,  -18'd6693,  -18'd2516,  18'd3131,  -18'd5100,  -18'd240,  -18'd9229,  -18'd1045,  
-18'd11579,  -18'd1008,  -18'd1300,  18'd27,  -18'd8521,  -18'd1515,  -18'd770,  -18'd13355,  -18'd6513,  -18'd5776,  18'd3867,  18'd4060,  -18'd6459,  18'd4623,  18'd5874,  -18'd5441,  
18'd3191,  18'd3772,  -18'd731,  -18'd80,  -18'd3041,  -18'd905,  -18'd8340,  -18'd5342,  18'd1106,  -18'd2777,  -18'd6249,  18'd2172,  18'd1313,  18'd4111,  -18'd5089,  18'd2343,  
18'd4334,  -18'd5237,  -18'd6924,  -18'd5691,  -18'd2071,  18'd6789,  18'd3256,  -18'd6481,  -18'd11205,  18'd4210,  -18'd4982,  18'd4048,  -18'd1772,  -18'd856,  -18'd10976,  -18'd10517,  
-18'd4736,  -18'd9743,  -18'd4682,  18'd6300,  -18'd6051,  -18'd5408,  -18'd1383,  18'd4433,  -18'd3242,  18'd5326,  -18'd6756,  18'd1282,  -18'd8068,  18'd11876,  -18'd6444,  18'd3219,  
-18'd9785,  -18'd5946,  -18'd9350,  18'd10061,  18'd7127,  18'd4395,  -18'd1666,  -18'd726,  -18'd2129,  -18'd1904,  18'd3202,  -18'd10968,  18'd455,  -18'd12143,  -18'd7725,  -18'd5664,  
18'd4741,  18'd1821,  -18'd10136,  18'd1417,  -18'd5473,  18'd3580,  -18'd8701,  18'd3752,  -18'd4212,  -18'd743,  -18'd6848,  18'd632,  18'd2664,  -18'd6958,  18'd4205,  -18'd7409,  
-18'd403,  18'd645,  18'd3874,  -18'd612,  18'd138,  18'd6000,  18'd5475,  18'd7491,  -18'd7377,  -18'd2865,  -18'd3497,  -18'd3274,  18'd1740,  18'd5293,  -18'd13205,  -18'd7106,  
18'd1803,  -18'd2657,  -18'd1150,  -18'd1644,  18'd5128,  -18'd2406,  -18'd8499,  -18'd6222,  -18'd5714,  18'd4655,  -18'd10289,  -18'd10635,  18'd3129,  -18'd6380,  18'd2491,  18'd7227,  

18'd3035,  18'd4759,  -18'd7139,  18'd2789,  18'd8166,  -18'd4511,  -18'd3360,  -18'd1141,  18'd648,  -18'd12597,  -18'd8154,  -18'd12826,  -18'd2338,  -18'd2690,  18'd3269,  -18'd9293,  
18'd5876,  -18'd9145,  -18'd10898,  18'd3123,  -18'd7135,  -18'd9288,  -18'd2493,  -18'd3029,  -18'd7050,  -18'd119,  18'd1065,  -18'd4436,  18'd7732,  18'd2821,  18'd3537,  -18'd5785,  
-18'd3765,  -18'd6955,  -18'd3794,  -18'd3247,  18'd5667,  -18'd3914,  -18'd2820,  18'd1567,  -18'd7982,  -18'd10930,  18'd5289,  -18'd4112,  18'd4529,  18'd6304,  18'd6675,  -18'd7184,  
18'd2233,  18'd3835,  -18'd4819,  -18'd2195,  -18'd2419,  18'd1122,  -18'd4235,  18'd3534,  -18'd9104,  -18'd4001,  18'd68,  18'd376,  -18'd3555,  -18'd2268,  18'd1763,  -18'd2788,  
-18'd12153,  -18'd8735,  18'd3486,  -18'd9168,  18'd5615,  -18'd6289,  -18'd2912,  18'd3836,  -18'd1815,  18'd1534,  -18'd6639,  -18'd746,  -18'd983,  -18'd612,  18'd680,  -18'd4177,  
-18'd3607,  -18'd7464,  18'd110,  18'd1032,  -18'd6718,  -18'd2401,  -18'd5979,  18'd4049,  18'd1027,  18'd4406,  -18'd9641,  -18'd1905,  18'd8473,  -18'd1205,  -18'd11426,  -18'd3178,  
18'd2798,  -18'd4310,  -18'd6466,  -18'd9983,  18'd1893,  18'd7659,  -18'd1663,  -18'd2918,  -18'd5708,  -18'd5748,  -18'd7916,  18'd1999,  18'd3465,  -18'd6701,  -18'd7687,  -18'd4910,  
-18'd10084,  18'd982,  18'd3054,  -18'd91,  18'd4173,  -18'd1970,  -18'd984,  -18'd7568,  18'd2005,  18'd4335,  18'd6305,  18'd1223,  -18'd4298,  -18'd11798,  -18'd4548,  18'd285,  
18'd2004,  -18'd9904,  -18'd4521,  -18'd518,  18'd4342,  -18'd8048,  -18'd1877,  -18'd8064,  18'd3769,  -18'd1922,  18'd2240,  18'd2974,  -18'd1808,  -18'd10234,  18'd1877,  -18'd3095,  
18'd4829,  18'd7916,  -18'd7116,  -18'd10550,  18'd6544,  -18'd463,  -18'd2455,  -18'd386,  18'd3011,  -18'd10581,  -18'd4101,  -18'd1060,  -18'd6230,  18'd3730,  18'd4111,  18'd1054,  
18'd1873,  -18'd3091,  18'd3750,  -18'd4084,  -18'd4725,  18'd4196,  -18'd12044,  -18'd9107,  -18'd4817,  -18'd3485,  -18'd2172,  18'd7435,  18'd8715,  18'd5351,  -18'd10776,  -18'd4164,  
18'd1307,  18'd649,  18'd5153,  -18'd4671,  18'd4198,  -18'd9865,  18'd1174,  18'd3612,  -18'd3757,  -18'd6836,  -18'd10218,  -18'd443,  18'd8936,  -18'd9890,  -18'd4429,  18'd5099,  
-18'd7816,  -18'd2104,  -18'd10316,  18'd58,  18'd5316,  -18'd7013,  -18'd3819,  18'd4969,  -18'd1505,  18'd400,  -18'd3246,  -18'd2583,  18'd6887,  18'd4925,  -18'd10563,  18'd6810,  
-18'd7002,  -18'd9125,  -18'd7162,  18'd5199,  -18'd2334,  -18'd7361,  -18'd10901,  -18'd7013,  -18'd4591,  -18'd1173,  -18'd10554,  -18'd4595,  -18'd1814,  -18'd2153,  -18'd6097,  -18'd2642,  
-18'd1548,  18'd3546,  18'd5139,  18'd4795,  18'd1958,  -18'd1565,  -18'd145,  -18'd2036,  -18'd4495,  18'd2679,  -18'd8931,  -18'd1846,  18'd2846,  18'd1307,  18'd3295,  -18'd7783,  
-18'd8504,  18'd4837,  18'd478,  -18'd7903,  -18'd4121,  -18'd10266,  18'd178,  -18'd8020,  -18'd9631,  -18'd6762,  -18'd1232,  18'd2047,  18'd6596,  -18'd2612,  18'd1647,  18'd5357,  

-18'd4893,  18'd18738,  18'd63,  -18'd20169,  18'd3514,  -18'd7683,  -18'd13233,  18'd6627,  -18'd17438,  18'd6602,  18'd8800,  18'd3422,  18'd2682,  -18'd9530,  18'd5792,  -18'd16623,  
-18'd3828,  -18'd94,  18'd7682,  -18'd29494,  -18'd3601,  -18'd6217,  -18'd4879,  18'd9679,  -18'd212,  -18'd11052,  -18'd2767,  -18'd7662,  18'd1295,  -18'd8016,  18'd3493,  -18'd2115,  
-18'd3317,  -18'd11386,  18'd2563,  -18'd25643,  -18'd2477,  -18'd1489,  -18'd5282,  18'd1260,  -18'd976,  18'd1654,  18'd2988,  -18'd10948,  -18'd2530,  18'd1261,  -18'd3436,  18'd8989,  
18'd2880,  -18'd3417,  18'd4701,  18'd1436,  -18'd4876,  18'd7866,  -18'd7727,  -18'd15034,  -18'd16369,  18'd26319,  18'd30209,  18'd10332,  -18'd5345,  -18'd7928,  18'd9979,  18'd9973,  
-18'd99,  18'd14844,  18'd3184,  -18'd20245,  -18'd5669,  -18'd4862,  18'd4019,  18'd7120,  18'd2076,  18'd22064,  18'd5622,  18'd10664,  -18'd6559,  -18'd2145,  18'd2414,  -18'd6015,  
18'd4952,  18'd5239,  -18'd1931,  -18'd12326,  18'd1225,  18'd117,  18'd2629,  -18'd4326,  -18'd8357,  -18'd16685,  -18'd12160,  -18'd12903,  -18'd8128,  18'd3686,  18'd1189,  -18'd7871,  
-18'd150,  -18'd5239,  18'd17457,  -18'd2117,  18'd4425,  -18'd9312,  18'd3503,  18'd15209,  18'd10265,  18'd4701,  -18'd5360,  -18'd621,  18'd5508,  -18'd5957,  18'd6450,  -18'd4392,  
18'd9971,  -18'd11472,  -18'd7122,  18'd7538,  18'd5238,  -18'd7108,  18'd26246,  -18'd8812,  18'd8576,  18'd1433,  18'd6361,  -18'd12015,  -18'd7359,  -18'd7143,  18'd12538,  -18'd2359,  
18'd988,  18'd4828,  18'd3536,  18'd7871,  18'd749,  -18'd322,  -18'd8752,  -18'd367,  18'd7757,  -18'd2045,  -18'd2205,  18'd3611,  -18'd7702,  18'd12187,  -18'd11532,  18'd8933,  
18'd9998,  -18'd693,  18'd3706,  18'd9975,  -18'd8494,  18'd2959,  18'd2467,  18'd7288,  18'd4474,  -18'd2078,  18'd3139,  18'd7023,  -18'd9408,  -18'd765,  -18'd4261,  18'd10057,  
-18'd2791,  18'd5969,  18'd2449,  18'd6046,  -18'd4213,  -18'd11684,  18'd1282,  18'd12011,  18'd7321,  -18'd2168,  18'd4557,  18'd5374,  18'd5705,  18'd5276,  18'd9401,  18'd13161,  
18'd1844,  18'd5890,  18'd1827,  18'd6711,  18'd5667,  18'd5307,  18'd13354,  18'd3983,  18'd2506,  -18'd884,  18'd3288,  -18'd5133,  -18'd4261,  -18'd9542,  -18'd3851,  -18'd2126,  
18'd8773,  18'd13471,  -18'd8796,  18'd20040,  -18'd5047,  18'd2886,  -18'd4301,  -18'd16454,  18'd14825,  18'd13999,  -18'd10150,  18'd13447,  -18'd2104,  18'd17680,  -18'd5006,  18'd10847,  
18'd1994,  18'd11503,  -18'd21753,  18'd11154,  18'd232,  -18'd9650,  -18'd20950,  18'd6759,  -18'd362,  18'd2626,  -18'd678,  18'd12940,  -18'd4246,  18'd19103,  -18'd10389,  18'd5003,  
-18'd11843,  18'd21149,  18'd1006,  18'd10965,  18'd2332,  -18'd2715,  18'd957,  18'd16056,  -18'd3339,  -18'd1879,  -18'd248,  -18'd2087,  18'd7845,  18'd2838,  -18'd6286,  18'd5016,  
-18'd11345,  18'd2881,  18'd6911,  18'd6723,  -18'd6958,  18'd5435,  -18'd2818,  18'd14655,  -18'd16142,  -18'd524,  18'd11673,  -18'd1871,  18'd3105,  18'd14992,  -18'd15836,  -18'd6687,  

18'd5127,  -18'd6477,  -18'd779,  -18'd5257,  -18'd2106,  18'd3991,  18'd2653,  18'd625,  -18'd6078,  -18'd3330,  -18'd3057,  -18'd3939,  18'd623,  -18'd6434,  -18'd8296,  -18'd9344,  
-18'd266,  -18'd4472,  -18'd5426,  18'd4118,  18'd1732,  18'd2715,  18'd301,  -18'd1166,  18'd2116,  18'd334,  18'd2223,  -18'd5745,  -18'd7811,  -18'd15,  -18'd83,  -18'd115,  
-18'd369,  18'd5494,  18'd274,  18'd3008,  18'd7532,  18'd3342,  -18'd9139,  -18'd9378,  18'd6181,  -18'd6678,  18'd2307,  18'd2582,  18'd1893,  18'd3342,  18'd6701,  -18'd8436,  
-18'd1440,  -18'd784,  18'd3558,  18'd6554,  -18'd2879,  18'd4622,  -18'd9847,  18'd1852,  18'd5141,  18'd1739,  18'd1464,  18'd5020,  18'd6152,  -18'd1875,  18'd7538,  18'd5691,  
-18'd8165,  -18'd4721,  -18'd9776,  -18'd1946,  -18'd7992,  -18'd6490,  18'd7120,  18'd756,  -18'd912,  -18'd5504,  -18'd3405,  18'd4138,  -18'd3488,  18'd283,  -18'd3014,  18'd5888,  
18'd234,  -18'd4486,  18'd2751,  18'd4766,  -18'd6830,  18'd450,  18'd4714,  -18'd7063,  -18'd3600,  18'd5376,  18'd3394,  -18'd6715,  18'd2861,  -18'd2775,  -18'd10106,  -18'd9703,  
-18'd2575,  18'd6436,  18'd5506,  -18'd9756,  -18'd2015,  18'd4835,  -18'd1483,  18'd5766,  -18'd934,  -18'd8883,  18'd2330,  18'd329,  -18'd7881,  18'd5819,  -18'd1325,  -18'd255,  
-18'd2996,  18'd7267,  -18'd4438,  18'd5512,  18'd8834,  -18'd8930,  -18'd4925,  -18'd151,  -18'd3086,  -18'd7778,  -18'd5924,  -18'd5938,  18'd7526,  -18'd6315,  18'd3252,  18'd2442,  
18'd5909,  18'd1164,  -18'd10025,  18'd1315,  18'd4204,  18'd6936,  18'd3666,  -18'd2817,  18'd2313,  -18'd10111,  -18'd7924,  -18'd8798,  -18'd7714,  18'd2250,  -18'd7931,  18'd2969,  
-18'd7202,  -18'd9289,  18'd6294,  18'd483,  18'd4256,  18'd3189,  -18'd8563,  18'd4466,  18'd5149,  18'd5380,  -18'd8928,  -18'd7575,  -18'd8636,  -18'd10381,  -18'd8672,  -18'd2861,  
-18'd10512,  -18'd8614,  18'd2419,  -18'd3401,  18'd2451,  -18'd8664,  -18'd8241,  -18'd4335,  -18'd4120,  -18'd7649,  18'd3579,  -18'd1647,  -18'd838,  18'd5727,  -18'd7337,  18'd5267,  
-18'd9579,  18'd2047,  -18'd6096,  -18'd543,  18'd4395,  -18'd6348,  18'd2825,  -18'd7550,  18'd2684,  -18'd2705,  -18'd2747,  18'd2840,  18'd5879,  -18'd6655,  -18'd10392,  -18'd651,  
-18'd3752,  -18'd9398,  18'd4192,  -18'd7183,  18'd2814,  -18'd4643,  -18'd4714,  18'd5589,  -18'd8763,  -18'd7892,  -18'd7220,  -18'd6921,  18'd7555,  -18'd511,  -18'd1184,  -18'd1875,  
-18'd4834,  -18'd3789,  -18'd7259,  18'd5448,  -18'd4131,  18'd614,  -18'd9402,  18'd4062,  -18'd7358,  -18'd8746,  18'd2921,  -18'd5014,  -18'd3435,  -18'd7264,  -18'd8472,  -18'd10687,  
18'd1210,  -18'd3093,  -18'd7741,  -18'd3793,  -18'd491,  18'd4967,  -18'd9711,  18'd348,  -18'd8630,  18'd7047,  -18'd2466,  18'd4427,  -18'd2711,  18'd4833,  18'd7224,  -18'd8076,  
-18'd6851,  -18'd4544,  18'd4740,  -18'd7001,  18'd7682,  -18'd2165,  18'd1411,  -18'd3790,  -18'd1233,  18'd4943,  18'd1282,  18'd5418,  -18'd3876,  -18'd1913,  18'd4955,  -18'd6611,  

-18'd1146,  -18'd5289,  -18'd4890,  18'd13333,  18'd1424,  18'd5039,  -18'd10943,  -18'd7769,  -18'd17791,  -18'd6216,  -18'd5949,  18'd489,  18'd1152,  18'd6338,  -18'd2726,  18'd27712,  
-18'd17544,  18'd20272,  -18'd2599,  -18'd1149,  18'd2289,  18'd719,  18'd2605,  18'd16706,  -18'd5428,  -18'd11783,  -18'd5399,  -18'd20902,  18'd4508,  -18'd4688,  18'd648,  18'd7453,  
18'd3404,  -18'd530,  -18'd776,  18'd14437,  18'd3919,  -18'd23791,  18'd4349,  -18'd256,  -18'd20688,  18'd10045,  18'd12072,  -18'd11453,  18'd5364,  -18'd17349,  18'd19720,  18'd4544,  
18'd6234,  -18'd12512,  -18'd15646,  18'd863,  18'd6560,  -18'd373,  18'd12512,  18'd749,  -18'd12692,  18'd8326,  18'd20933,  -18'd27324,  -18'd5005,  -18'd4362,  18'd16699,  -18'd192,  
-18'd4655,  18'd8269,  18'd4374,  18'd30753,  -18'd6085,  18'd3431,  18'd8730,  -18'd4666,  18'd7520,  18'd13942,  18'd10878,  -18'd5970,  -18'd3651,  18'd1850,  18'd5026,  -18'd13712,  
18'd4950,  18'd2279,  -18'd603,  18'd17586,  -18'd373,  18'd5501,  18'd8980,  18'd11663,  18'd18150,  18'd5640,  18'd12685,  18'd2394,  18'd1594,  -18'd3230,  18'd5891,  18'd2273,  
18'd4521,  18'd10122,  18'd9255,  18'd12132,  -18'd7573,  -18'd2161,  18'd13569,  18'd15211,  -18'd5252,  18'd1111,  18'd14209,  18'd7762,  18'd105,  18'd2191,  18'd5448,  -18'd2955,  
18'd15853,  -18'd7343,  18'd20505,  -18'd6053,  -18'd1579,  18'd11700,  18'd25815,  18'd7912,  18'd2623,  -18'd1233,  18'd25059,  18'd11477,  -18'd10333,  -18'd1437,  18'd10677,  18'd973,  
18'd5146,  -18'd4495,  18'd2353,  18'd9182,  -18'd5278,  -18'd620,  18'd11037,  18'd1214,  18'd9886,  18'd12328,  18'd6225,  18'd7844,  -18'd3325,  18'd4378,  -18'd1696,  -18'd17182,  
-18'd7084,  18'd3506,  18'd12569,  18'd2404,  -18'd7128,  18'd13142,  18'd24989,  -18'd11543,  18'd11498,  18'd6518,  18'd13403,  -18'd1374,  18'd3261,  -18'd6937,  18'd3598,  -18'd5318,  
-18'd6326,  -18'd4118,  18'd920,  -18'd655,  -18'd550,  -18'd3920,  18'd1289,  -18'd11453,  18'd6434,  -18'd8458,  -18'd2682,  18'd2486,  -18'd1404,  18'd5285,  -18'd3990,  18'd6066,  
18'd3314,  18'd908,  18'd1719,  18'd1064,  -18'd2633,  -18'd13557,  -18'd11831,  -18'd11923,  18'd4103,  -18'd2699,  18'd6189,  18'd4879,  18'd5509,  18'd1998,  -18'd9271,  -18'd6536,  
-18'd8537,  -18'd9283,  18'd4284,  -18'd5782,  18'd6842,  18'd9509,  18'd4672,  -18'd6657,  18'd5172,  -18'd10510,  -18'd8190,  -18'd5470,  -18'd3380,  18'd11234,  -18'd2146,  -18'd14987,  
-18'd395,  18'd13478,  18'd10257,  -18'd6878,  18'd389,  18'd25155,  18'd11561,  18'd4996,  18'd15981,  -18'd21658,  -18'd13706,  18'd3200,  -18'd3866,  18'd16744,  18'd824,  -18'd1472,  
-18'd1803,  18'd2051,  18'd2015,  18'd4450,  18'd8744,  18'd20726,  18'd13856,  -18'd8091,  -18'd817,  -18'd10793,  -18'd7263,  18'd689,  -18'd11082,  18'd16031,  -18'd14050,  18'd10592,  
18'd9078,  18'd4843,  -18'd10856,  18'd5386,  -18'd514,  18'd11240,  -18'd6488,  -18'd5634,  18'd7998,  18'd8028,  18'd3628,  -18'd4980,  18'd6167,  18'd5880,  -18'd7820,  18'd10270,  

18'd10919,  -18'd23392,  -18'd13730,  -18'd1701,  18'd8275,  -18'd4470,  -18'd10698,  18'd2216,  -18'd5243,  18'd20478,  -18'd3680,  18'd14056,  18'd4593,  18'd22538,  -18'd234,  -18'd20407,  
18'd5409,  -18'd13794,  -18'd4037,  18'd12332,  18'd9048,  -18'd2478,  18'd3834,  18'd7405,  -18'd8377,  -18'd44,  -18'd3189,  -18'd2020,  -18'd1408,  -18'd1129,  18'd1118,  -18'd1291,  
-18'd5724,  -18'd19910,  -18'd2036,  -18'd3356,  18'd9069,  -18'd15084,  18'd3010,  18'd10092,  18'd1875,  18'd16071,  18'd11175,  18'd7932,  -18'd1814,  -18'd15801,  18'd28420,  18'd345,  
18'd4786,  -18'd15173,  -18'd354,  -18'd6498,  18'd7602,  -18'd8139,  18'd1892,  18'd13235,  18'd13422,  18'd5258,  18'd29047,  18'd28505,  -18'd4577,  -18'd1121,  18'd27893,  -18'd13441,  
-18'd5674,  -18'd2888,  -18'd10304,  -18'd3044,  -18'd4460,  18'd4202,  -18'd1581,  18'd696,  -18'd1488,  18'd15693,  -18'd6207,  18'd13092,  18'd2761,  -18'd1865,  18'd10137,  -18'd14677,  
18'd1169,  18'd4641,  -18'd1288,  18'd1204,  18'd3350,  -18'd8817,  18'd2867,  18'd3325,  -18'd8102,  18'd7005,  -18'd1225,  -18'd3110,  -18'd1221,  -18'd12600,  18'd1465,  -18'd4650,  
18'd3473,  18'd1701,  18'd10968,  18'd970,  18'd2733,  -18'd12646,  -18'd9918,  18'd11804,  18'd551,  18'd3294,  18'd1380,  18'd17786,  -18'd2383,  -18'd11640,  18'd5730,  -18'd11234,  
18'd5769,  18'd8716,  18'd20837,  -18'd10665,  18'd6510,  -18'd15242,  18'd10171,  18'd17682,  -18'd7983,  18'd5297,  18'd3397,  18'd16818,  -18'd1728,  -18'd10907,  18'd11923,  18'd10442,  
-18'd10137,  18'd12527,  18'd9110,  -18'd16698,  18'd966,  -18'd8483,  -18'd364,  -18'd2246,  -18'd7050,  -18'd7833,  18'd11988,  18'd7097,  18'd3310,  18'd10803,  -18'd1325,  -18'd9824,  
18'd2730,  18'd6353,  18'd6940,  18'd8400,  18'd1759,  18'd19116,  18'd10299,  -18'd8655,  -18'd1534,  -18'd4191,  -18'd5687,  18'd1744,  18'd3777,  18'd10293,  -18'd13689,  -18'd10984,  
18'd9600,  18'd5402,  -18'd6729,  -18'd1631,  18'd4300,  -18'd1253,  18'd4128,  -18'd4309,  18'd8320,  18'd5338,  -18'd7907,  18'd3440,  -18'd1052,  18'd6427,  18'd3276,  -18'd2898,  
-18'd1288,  -18'd3898,  18'd24283,  -18'd12708,  -18'd8526,  -18'd14343,  -18'd10496,  18'd12219,  -18'd19500,  -18'd3500,  -18'd4731,  18'd270,  -18'd1361,  -18'd296,  -18'd10141,  -18'd8898,  
-18'd11837,  18'd2172,  18'd8035,  18'd4819,  -18'd736,  -18'd2821,  18'd605,  18'd7213,  18'd1730,  -18'd268,  18'd4906,  18'd4349,  18'd8455,  18'd12800,  18'd8675,  18'd14334,  
18'd6911,  18'd2664,  -18'd2733,  18'd1316,  18'd8228,  18'd10748,  -18'd11042,  -18'd1257,  18'd1122,  -18'd4037,  -18'd3851,  18'd8459,  18'd1192,  18'd13835,  -18'd966,  18'd13085,  
18'd5542,  18'd1565,  18'd6927,  18'd4317,  -18'd6396,  18'd10293,  18'd4528,  18'd9720,  18'd6834,  18'd301,  18'd3354,  -18'd8259,  -18'd6332,  18'd7770,  -18'd4840,  -18'd243,  
18'd2609,  18'd13792,  18'd3859,  -18'd8783,  18'd4606,  -18'd10195,  18'd936,  -18'd2899,  -18'd6791,  18'd6163,  -18'd1477,  18'd5358,  -18'd3301,  18'd13413,  18'd4237,  18'd15260,  

-18'd2789,  -18'd7174,  18'd2042,  -18'd17019,  -18'd1042,  -18'd1869,  18'd6664,  -18'd3066,  -18'd9139,  18'd16315,  18'd8646,  18'd3834,  18'd4162,  18'd3307,  18'd7469,  -18'd33601,  
18'd8320,  -18'd6634,  18'd220,  18'd6031,  18'd3494,  -18'd2579,  18'd4245,  -18'd14577,  18'd15252,  18'd11615,  -18'd2933,  18'd14074,  -18'd22,  -18'd8715,  18'd8949,  -18'd11686,  
18'd10046,  -18'd9017,  18'd6797,  18'd1119,  18'd4525,  18'd13752,  18'd9335,  -18'd11309,  18'd7136,  18'd8819,  18'd3488,  18'd16044,  -18'd894,  -18'd1138,  18'd5639,  18'd1982,  
18'd17241,  -18'd19692,  18'd6484,  -18'd4936,  18'd631,  18'd6647,  18'd1131,  -18'd8870,  18'd12189,  -18'd5367,  18'd18821,  18'd31606,  -18'd4061,  18'd5350,  18'd19099,  18'd2461,  
-18'd14850,  18'd7515,  18'd4367,  -18'd26557,  18'd2975,  -18'd6641,  18'd3879,  -18'd2222,  -18'd1767,  18'd8813,  18'd4238,  -18'd1434,  18'd2200,  -18'd9773,  18'd2894,  -18'd3084,  
-18'd7800,  18'd5059,  18'd9132,  -18'd5328,  18'd2171,  -18'd6255,  18'd239,  18'd3038,  -18'd7382,  18'd23389,  18'd3529,  -18'd5785,  18'd1458,  18'd4358,  18'd3203,  -18'd5933,  
-18'd1870,  -18'd12309,  18'd5477,  -18'd1017,  18'd7438,  -18'd2424,  18'd9373,  -18'd105,  18'd13441,  -18'd5122,  18'd9420,  -18'd5318,  -18'd6311,  -18'd6990,  18'd3886,  -18'd6286,  
18'd9287,  -18'd1064,  18'd20744,  -18'd1011,  18'd7346,  -18'd8831,  18'd5421,  18'd507,  18'd8154,  -18'd21896,  18'd4123,  -18'd8475,  -18'd178,  -18'd10100,  18'd15193,  18'd16627,  
-18'd8604,  18'd19059,  -18'd1258,  -18'd7992,  18'd4821,  -18'd7250,  18'd6488,  18'd11548,  18'd765,  18'd8873,  -18'd1725,  18'd5534,  18'd4349,  18'd11801,  18'd5149,  18'd6901,  
-18'd7982,  18'd4578,  18'd7549,  -18'd5944,  -18'd5398,  18'd6410,  -18'd14339,  -18'd1630,  18'd2376,  18'd4325,  18'd5753,  18'd18149,  18'd9584,  18'd6429,  -18'd4978,  18'd4609,  
18'd4735,  18'd2565,  18'd7,  -18'd5100,  -18'd2400,  18'd3003,  -18'd18086,  18'd15615,  -18'd7665,  18'd840,  -18'd2057,  18'd1715,  18'd3937,  18'd2507,  -18'd4755,  -18'd14679,  
18'd597,  18'd8065,  18'd20546,  18'd9714,  18'd5,  -18'd3490,  18'd7120,  18'd24107,  18'd6255,  -18'd27553,  18'd8950,  -18'd13346,  -18'd7641,  18'd2015,  -18'd870,  -18'd7765,  
18'd2581,  -18'd7601,  -18'd2874,  -18'd3983,  -18'd8416,  -18'd3357,  18'd2409,  18'd6755,  18'd1466,  -18'd8701,  -18'd534,  -18'd3822,  18'd6673,  -18'd1948,  18'd5417,  18'd3386,  
18'd44,  18'd6673,  -18'd9271,  -18'd8347,  -18'd7537,  18'd5335,  -18'd7596,  18'd383,  -18'd1169,  18'd16753,  -18'd4735,  18'd490,  18'd2256,  18'd11776,  -18'd6226,  18'd2696,  
-18'd953,  -18'd2966,  -18'd26436,  18'd14402,  -18'd5650,  -18'd4582,  -18'd24157,  18'd3824,  18'd5207,  18'd1892,  -18'd8057,  -18'd10014,  18'd2693,  18'd2822,  18'd6130,  18'd2737,  
-18'd4598,  18'd14690,  -18'd13128,  18'd2383,  18'd3758,  18'd14715,  18'd2295,  -18'd1738,  18'd963,  -18'd21794,  -18'd4338,  -18'd4535,  18'd7339,  -18'd2155,  -18'd11299,  -18'd4192,  

-18'd30961,  -18'd10357,  18'd5180,  -18'd7678,  -18'd6440,  -18'd13082,  18'd3489,  18'd1532,  -18'd27947,  -18'd12247,  18'd12862,  -18'd28796,  -18'd4504,  -18'd30961,  18'd4957,  -18'd4561,  
-18'd20718,  18'd16111,  18'd1719,  -18'd32415,  -18'd7116,  18'd6148,  18'd22865,  18'd11051,  18'd13649,  -18'd2148,  18'd2900,  18'd153,  18'd4107,  -18'd6458,  -18'd7173,  18'd3218,  
18'd8333,  18'd9081,  -18'd8393,  -18'd12302,  18'd1141,  18'd28608,  18'd14523,  -18'd16738,  18'd19737,  18'd9425,  -18'd2516,  18'd238,  -18'd4085,  18'd3375,  -18'd9327,  -18'd10179,  
18'd20005,  -18'd7055,  -18'd739,  -18'd10567,  -18'd7856,  18'd8994,  -18'd11804,  -18'd18000,  18'd2580,  -18'd529,  18'd7594,  -18'd2707,  18'd4316,  18'd5380,  18'd6565,  18'd7964,  
-18'd28312,  18'd1697,  18'd11228,  18'd24,  -18'd4762,  18'd8030,  18'd1023,  -18'd2720,  18'd17916,  -18'd365,  18'd9070,  18'd13360,  18'd4764,  18'd1825,  -18'd3245,  18'd1084,  
-18'd5276,  18'd743,  18'd812,  -18'd3617,  -18'd4418,  -18'd4157,  -18'd9057,  18'd12042,  -18'd10405,  -18'd8224,  -18'd9772,  -18'd13026,  -18'd2901,  18'd5684,  18'd6006,  18'd9804,  
-18'd8540,  18'd14041,  -18'd1923,  -18'd4346,  18'd9197,  18'd24043,  -18'd4398,  18'd427,  18'd935,  18'd11651,  18'd5645,  18'd350,  18'd8063,  18'd7965,  -18'd4113,  18'd7707,  
18'd12737,  18'd7356,  18'd7496,  18'd8406,  -18'd2337,  18'd8768,  18'd4617,  18'd14997,  18'd20069,  -18'd25683,  18'd3468,  18'd4124,  -18'd5576,  18'd7132,  -18'd4692,  18'd88,  
-18'd12697,  -18'd4068,  -18'd934,  18'd5549,  -18'd3522,  18'd4170,  18'd5909,  18'd74,  18'd2337,  -18'd1803,  -18'd5589,  18'd5865,  -18'd578,  -18'd3657,  18'd3062,  -18'd3339,  
18'd7814,  -18'd3087,  -18'd3254,  18'd6127,  18'd3209,  -18'd3072,  -18'd15892,  -18'd14128,  -18'd13670,  -18'd4055,  -18'd5109,  -18'd10503,  -18'd6907,  -18'd1181,  18'd851,  18'd2447,  
18'd3847,  18'd17852,  -18'd2882,  -18'd464,  18'd4443,  -18'd786,  -18'd6328,  18'd15520,  18'd834,  -18'd350,  -18'd3357,  18'd6187,  -18'd7672,  18'd15308,  18'd6188,  18'd723,  
18'd4428,  18'd7760,  18'd9936,  18'd12619,  -18'd4956,  18'd8774,  -18'd1728,  18'd6450,  18'd8184,  -18'd5526,  18'd13936,  -18'd2672,  -18'd402,  -18'd8928,  18'd13886,  18'd13145,  
18'd754,  -18'd11682,  -18'd2118,  -18'd24504,  18'd1024,  18'd12847,  18'd5905,  -18'd4333,  18'd618,  18'd3818,  -18'd1143,  -18'd1019,  18'd322,  -18'd8655,  18'd7136,  -18'd11638,  
18'd679,  -18'd3890,  18'd1514,  -18'd13040,  -18'd8192,  -18'd3385,  -18'd5938,  -18'd423,  -18'd10965,  -18'd734,  18'd4787,  -18'd15757,  18'd5582,  -18'd962,  18'd7393,  18'd6254,  
18'd15671,  -18'd1490,  -18'd17568,  -18'd10501,  18'd3615,  -18'd21089,  -18'd12459,  -18'd1865,  -18'd6145,  18'd3435,  -18'd84,  18'd10934,  18'd2641,  18'd2043,  18'd14422,  18'd1249,  
18'd7344,  18'd9255,  18'd4404,  18'd8634,  18'd8956,  -18'd4390,  18'd2922,  18'd4535,  18'd21520,  -18'd3801,  18'd5414,  -18'd4356,  -18'd3267,  -18'd3010,  -18'd5477,  18'd4917,  

18'd23528,  18'd1181,  -18'd12940,  -18'd18327,  -18'd3468,  18'd7931,  -18'd10571,  -18'd1235,  18'd10725,  18'd6238,  -18'd4208,  18'd27397,  -18'd3922,  18'd14395,  -18'd13854,  18'd20469,  
18'd15285,  -18'd4540,  -18'd10734,  -18'd7328,  18'd2652,  -18'd8422,  -18'd13664,  -18'd15654,  18'd4872,  -18'd175,  -18'd10195,  18'd15029,  18'd73,  18'd19404,  -18'd16217,  18'd18223,  
18'd10903,  -18'd18879,  18'd6586,  18'd7074,  18'd1133,  -18'd15060,  -18'd10037,  -18'd27530,  18'd367,  18'd9431,  -18'd1400,  18'd11325,  -18'd815,  18'd8827,  -18'd12807,  18'd10359,  
-18'd4353,  -18'd9850,  18'd5008,  18'd11771,  18'd2734,  18'd4281,  -18'd8414,  -18'd18588,  18'd14242,  18'd12024,  18'd16685,  -18'd6758,  -18'd596,  18'd4560,  -18'd17655,  18'd15949,  
18'd19949,  -18'd12632,  -18'd7647,  -18'd731,  -18'd8558,  18'd7953,  18'd11542,  -18'd11377,  18'd10824,  18'd15186,  18'd3641,  -18'd3286,  18'd1262,  -18'd6636,  18'd6556,  -18'd12023,  
18'd8825,  -18'd4408,  -18'd12037,  18'd18536,  18'd3645,  -18'd4305,  -18'd2683,  18'd2545,  18'd14229,  -18'd10841,  -18'd3192,  -18'd4010,  -18'd4478,  -18'd7696,  18'd2695,  -18'd123,  
-18'd4461,  -18'd15374,  -18'd146,  18'd3414,  -18'd4211,  -18'd11825,  18'd5167,  -18'd7595,  18'd207,  18'd30010,  18'd3311,  18'd4979,  18'd3971,  -18'd12799,  -18'd3380,  -18'd2880,  
-18'd11332,  -18'd8008,  -18'd12281,  -18'd11037,  -18'd4554,  18'd4002,  -18'd6015,  -18'd14789,  -18'd2678,  18'd8976,  18'd19934,  18'd4732,  -18'd3616,  -18'd3143,  -18'd4016,  -18'd15752,  
-18'd6899,  -18'd1735,  18'd9668,  18'd7269,  -18'd7830,  18'd12608,  18'd24199,  -18'd3048,  18'd5077,  18'd11575,  18'd7158,  18'd11205,  -18'd6564,  18'd98,  18'd10285,  -18'd8043,  
18'd5604,  -18'd3030,  -18'd129,  18'd8072,  18'd7597,  -18'd681,  18'd21389,  -18'd3122,  18'd17873,  -18'd4006,  18'd14015,  -18'd14733,  18'd4879,  -18'd15802,  18'd5331,  18'd11240,  
-18'd4633,  -18'd15604,  18'd268,  -18'd3574,  -18'd5872,  -18'd11886,  18'd12195,  -18'd14510,  18'd442,  -18'd11722,  18'd7105,  -18'd16591,  18'd2092,  -18'd7773,  -18'd10687,  -18'd4546,  
18'd3446,  -18'd6661,  -18'd3364,  -18'd9113,  18'd2210,  -18'd8179,  -18'd3659,  -18'd12143,  -18'd587,  18'd167,  18'd7659,  18'd9191,  -18'd8537,  18'd540,  18'd9977,  -18'd12534,  
-18'd1912,  18'd3031,  18'd3676,  18'd14269,  18'd4262,  18'd7282,  18'd10569,  18'd4514,  18'd8890,  18'd8181,  18'd3109,  18'd25521,  -18'd9029,  -18'd11383,  -18'd58,  -18'd5248,  
-18'd4246,  -18'd1152,  18'd4568,  -18'd7955,  18'd120,  18'd6325,  18'd7195,  18'd8213,  18'd10410,  -18'd5208,  18'd10415,  18'd9711,  -18'd9493,  18'd5274,  18'd5148,  18'd4158,  
-18'd826,  -18'd5090,  -18'd3457,  -18'd4488,  -18'd6407,  18'd26241,  18'd19419,  -18'd181,  18'd5929,  -18'd10919,  18'd5043,  -18'd5808,  18'd5161,  18'd3639,  -18'd10578,  18'd426,  
18'd11138,  -18'd12855,  18'd2404,  -18'd13367,  18'd5489,  18'd19474,  18'd8951,  18'd4688,  18'd13871,  18'd4605,  -18'd5997,  18'd6784,  -18'd6217,  18'd1925,  -18'd1587,  -18'd2275,  

-18'd8998,  18'd16413,  18'd16964,  -18'd11760,  -18'd2694,  18'd20142,  18'd15276,  18'd11762,  18'd4551,  18'd6508,  18'd18495,  18'd11015,  18'd1227,  18'd1502,  18'd1963,  18'd20613,  
-18'd1151,  18'd10483,  18'd18808,  -18'd16588,  -18'd2,  18'd7015,  18'd9010,  18'd7805,  18'd30485,  -18'd748,  18'd6718,  -18'd6275,  -18'd10700,  18'd16997,  -18'd11942,  18'd34717,  
-18'd949,  18'd6041,  18'd89,  18'd14793,  -18'd7410,  18'd7420,  18'd1598,  -18'd19728,  18'd16242,  18'd9837,  18'd21765,  -18'd5866,  18'd5049,  18'd14771,  -18'd733,  18'd20325,  
18'd490,  -18'd12143,  -18'd2619,  18'd13574,  18'd1167,  -18'd4064,  -18'd16014,  -18'd46632,  18'd2380,  18'd21192,  18'd19723,  -18'd5658,  18'd3717,  -18'd1893,  18'd8689,  18'd10691,  
-18'd1224,  18'd8922,  18'd1803,  -18'd10634,  18'd918,  18'd9698,  -18'd249,  18'd4697,  18'd12890,  18'd5346,  18'd1153,  18'd3889,  -18'd5036,  18'd10612,  -18'd4676,  18'd6047,  
-18'd7992,  18'd962,  -18'd4860,  -18'd4951,  18'd1765,  18'd14882,  -18'd6557,  18'd10790,  18'd20060,  -18'd1580,  18'd19801,  18'd13488,  -18'd2627,  18'd7307,  18'd5037,  18'd9966,  
18'd4178,  -18'd7400,  18'd15256,  -18'd5237,  -18'd5390,  -18'd409,  18'd7986,  -18'd3289,  18'd29328,  -18'd8846,  18'd21627,  -18'd10721,  18'd6629,  -18'd1911,  18'd156,  -18'd4365,  
18'd7424,  18'd6972,  18'd5485,  18'd1459,  18'd8398,  18'd4756,  18'd1852,  -18'd2819,  -18'd814,  -18'd12145,  18'd6145,  -18'd6825,  -18'd433,  18'd1581,  18'd568,  -18'd2603,  
18'd7233,  18'd14004,  18'd486,  18'd19690,  18'd1204,  18'd5144,  -18'd11474,  18'd1872,  -18'd2858,  18'd694,  -18'd4952,  18'd9650,  18'd1820,  -18'd3754,  18'd2537,  18'd9630,  
18'd13831,  18'd7452,  -18'd356,  18'd4011,  18'd4439,  18'd2188,  18'd2194,  18'd1632,  -18'd8358,  18'd9077,  18'd2522,  18'd1407,  -18'd8894,  18'd183,  -18'd5079,  18'd4034,  
-18'd14079,  -18'd4322,  18'd9329,  18'd3287,  18'd4747,  18'd15,  18'd1211,  18'd3945,  18'd2449,  -18'd14804,  18'd613,  -18'd12674,  -18'd9413,  -18'd102,  18'd9068,  18'd6570,  
-18'd1801,  18'd26639,  18'd1364,  -18'd395,  18'd178,  -18'd15591,  -18'd10703,  18'd15493,  18'd7877,  -18'd10643,  -18'd11593,  18'd3210,  -18'd2577,  -18'd14625,  -18'd2991,  18'd6670,  
-18'd4077,  -18'd2799,  -18'd12527,  18'd7737,  18'd6515,  -18'd6156,  -18'd21389,  -18'd13587,  18'd6701,  -18'd2724,  -18'd19013,  -18'd3901,  -18'd2466,  18'd7490,  -18'd11621,  18'd1285,  
18'd2841,  18'd1519,  -18'd23486,  18'd1772,  18'd7294,  -18'd13938,  -18'd7256,  -18'd6385,  -18'd8561,  18'd1664,  -18'd9999,  18'd2669,  -18'd1732,  -18'd10341,  18'd11216,  -18'd1520,  
-18'd22873,  -18'd2056,  -18'd7102,  -18'd20663,  18'd807,  -18'd19063,  -18'd229,  18'd20182,  -18'd3094,  18'd4692,  -18'd5772,  -18'd4221,  -18'd4623,  -18'd7455,  -18'd7604,  -18'd19463,  
-18'd24040,  -18'd6550,  -18'd12815,  18'd10041,  -18'd5981,  -18'd19714,  -18'd12666,  18'd16288,  -18'd11290,  18'd5196,  -18'd7399,  -18'd8263,  18'd6780,  -18'd7310,  18'd2089,  -18'd2326,  

18'd8332,  -18'd11796,  -18'd8313,  -18'd25322,  -18'd1523,  -18'd2113,  18'd4129,  18'd8052,  -18'd10323,  18'd8210,  18'd13764,  18'd18198,  18'd8145,  -18'd20241,  18'd8882,  -18'd43959,  
-18'd4288,  -18'd18853,  18'd7616,  -18'd15308,  -18'd1923,  18'd18243,  18'd6694,  -18'd7095,  18'd32347,  18'd17091,  18'd11868,  18'd10241,  18'd2286,  -18'd2634,  18'd8507,  -18'd18913,  
18'd5628,  -18'd19424,  -18'd11783,  18'd11578,  -18'd2216,  -18'd4619,  -18'd11118,  -18'd11779,  18'd18464,  18'd15468,  18'd583,  18'd8513,  -18'd797,  -18'd2936,  18'd2286,  18'd3061,  
18'd11931,  -18'd8760,  -18'd1143,  18'd22707,  18'd4136,  -18'd2669,  -18'd5486,  -18'd2855,  18'd8773,  18'd21729,  18'd8933,  18'd10832,  -18'd2029,  18'd7945,  -18'd6369,  18'd5837,  
-18'd14057,  18'd11391,  18'd29,  -18'd31124,  -18'd7697,  -18'd9143,  -18'd3589,  18'd12079,  -18'd15700,  -18'd24092,  18'd6226,  -18'd6937,  18'd348,  -18'd26756,  -18'd1091,  18'd3187,  
-18'd15878,  -18'd1574,  18'd8976,  -18'd49897,  18'd3356,  -18'd3163,  18'd9433,  -18'd387,  18'd5338,  -18'd13972,  18'd4901,  -18'd14130,  -18'd6384,  18'd348,  18'd15605,  -18'd16847,  
-18'd3857,  -18'd6573,  18'd12936,  -18'd11242,  18'd4565,  -18'd1629,  -18'd2603,  -18'd2088,  18'd12695,  18'd19784,  -18'd1629,  18'd2519,  18'd9675,  -18'd12184,  18'd173,  -18'd8773,  
18'd9683,  18'd1662,  -18'd22826,  18'd19282,  -18'd1254,  -18'd2239,  -18'd7588,  18'd1547,  18'd10267,  18'd3500,  -18'd8169,  -18'd5142,  18'd6528,  -18'd2876,  -18'd2272,  -18'd10807,  
-18'd10191,  18'd2801,  18'd1892,  18'd8317,  -18'd301,  18'd628,  18'd10357,  18'd6325,  -18'd1669,  -18'd15550,  18'd211,  -18'd6995,  18'd7131,  -18'd12581,  -18'd1066,  18'd356,  
-18'd321,  18'd6335,  -18'd1581,  -18'd9289,  18'd989,  18'd56,  18'd6134,  -18'd17910,  -18'd6318,  18'd9361,  -18'd7176,  18'd8605,  -18'd7446,  -18'd12720,  18'd5880,  18'd2864,  
18'd8902,  18'd6318,  18'd6102,  -18'd6571,  18'd5394,  -18'd3289,  18'd15787,  -18'd9748,  18'd2325,  18'd6172,  -18'd5558,  -18'd3011,  -18'd116,  18'd8246,  -18'd666,  -18'd2121,  
-18'd98,  -18'd6123,  18'd9452,  18'd1767,  -18'd4254,  18'd352,  18'd16020,  -18'd5518,  18'd21699,  -18'd53,  -18'd687,  -18'd20562,  -18'd1423,  18'd1367,  18'd11688,  -18'd6119,  
18'd10131,  18'd3794,  18'd13605,  18'd13749,  18'd1439,  18'd18212,  -18'd5664,  -18'd8349,  18'd6696,  -18'd255,  -18'd375,  18'd11760,  18'd1989,  -18'd6600,  18'd1391,  18'd10458,  
-18'd1669,  18'd13448,  18'd9016,  -18'd10238,  -18'd6733,  18'd13359,  -18'd4070,  -18'd12162,  18'd422,  18'd14963,  18'd6256,  18'd14984,  18'd744,  -18'd5695,  -18'd5219,  18'd5584,  
18'd16068,  18'd3594,  -18'd9157,  -18'd3459,  -18'd6463,  18'd7320,  18'd11682,  18'd6218,  18'd8457,  -18'd314,  18'd8391,  18'd4023,  18'd8111,  18'd8312,  18'd6835,  18'd11590,  
-18'd5217,  18'd16273,  18'd22011,  -18'd5368,  18'd4825,  18'd4987,  18'd21864,  -18'd8293,  -18'd3877,  -18'd1555,  -18'd1542,  18'd4078,  18'd6738,  -18'd2018,  -18'd6459,  18'd1547,  

-18'd1065,  -18'd2885,  18'd4615,  18'd5382,  -18'd484,  18'd3584,  18'd2755,  -18'd10342,  18'd3490,  -18'd2784,  -18'd2220,  18'd6211,  18'd6930,  18'd2198,  -18'd3223,  18'd5780,  
18'd1323,  18'd1177,  -18'd6178,  -18'd7686,  18'd2506,  18'd3021,  -18'd6175,  -18'd8967,  18'd5727,  -18'd6296,  18'd3475,  18'd323,  -18'd2486,  18'd8459,  18'd3778,  18'd8539,  
-18'd6609,  -18'd5397,  -18'd3271,  18'd5694,  18'd6293,  18'd7274,  -18'd8890,  -18'd9069,  18'd161,  18'd2244,  -18'd5959,  -18'd9729,  -18'd2549,  -18'd5549,  18'd679,  -18'd8660,  
-18'd1392,  18'd933,  18'd4725,  -18'd1815,  18'd1867,  18'd2398,  18'd6477,  -18'd3092,  -18'd5339,  -18'd3053,  18'd4276,  18'd152,  -18'd4449,  -18'd7356,  -18'd1836,  18'd2773,  
18'd2692,  -18'd8986,  -18'd10451,  -18'd8068,  18'd8139,  -18'd5082,  -18'd4594,  18'd6177,  18'd6848,  -18'd7749,  -18'd6977,  -18'd3197,  18'd6117,  18'd4443,  18'd3071,  -18'd2999,  
-18'd3203,  -18'd6243,  -18'd1732,  -18'd3745,  18'd8340,  18'd4455,  -18'd2567,  18'd595,  -18'd5064,  18'd126,  -18'd2168,  -18'd5255,  -18'd1425,  -18'd3488,  -18'd8110,  -18'd716,  
-18'd7458,  -18'd8083,  -18'd10915,  18'd1910,  -18'd7425,  -18'd1629,  -18'd8851,  -18'd2424,  -18'd2833,  -18'd2120,  -18'd8629,  18'd2485,  18'd8960,  -18'd6351,  -18'd5406,  18'd3533,  
18'd4987,  18'd3454,  -18'd7464,  18'd240,  -18'd6879,  18'd5834,  -18'd8003,  -18'd1703,  18'd746,  -18'd6857,  -18'd2259,  -18'd6539,  18'd4453,  -18'd7297,  18'd4944,  -18'd7151,  
18'd2693,  -18'd3172,  -18'd3805,  -18'd3264,  18'd4545,  18'd2255,  -18'd4921,  -18'd8008,  -18'd2593,  -18'd2453,  -18'd9193,  18'd7029,  18'd1881,  -18'd6567,  -18'd4441,  -18'd4418,  
-18'd2522,  -18'd3894,  -18'd6984,  -18'd1781,  -18'd4282,  -18'd1312,  18'd6205,  -18'd6556,  18'd6314,  -18'd2547,  -18'd8222,  -18'd10306,  18'd1655,  18'd4860,  -18'd2039,  -18'd5361,  
18'd5318,  -18'd3750,  -18'd9461,  18'd5538,  18'd6098,  18'd3273,  18'd3404,  -18'd1650,  -18'd1009,  18'd1404,  18'd2543,  18'd453,  -18'd8166,  18'd7861,  18'd3329,  -18'd8926,  
18'd6947,  -18'd1101,  -18'd7029,  -18'd7143,  18'd1211,  18'd8797,  18'd2663,  -18'd5393,  18'd4211,  -18'd9711,  -18'd9083,  18'd6621,  -18'd8816,  18'd656,  18'd6429,  -18'd695,  
18'd36,  -18'd4581,  18'd6081,  18'd1633,  18'd432,  -18'd4350,  -18'd3553,  -18'd3710,  -18'd1267,  -18'd6079,  -18'd4855,  18'd5744,  18'd2808,  -18'd9063,  18'd3511,  -18'd2545,  
-18'd2100,  -18'd5854,  18'd4649,  18'd6444,  -18'd3941,  -18'd8628,  -18'd1726,  -18'd11031,  18'd194,  -18'd7419,  18'd5828,  -18'd5248,  -18'd5384,  -18'd480,  -18'd2428,  18'd3397,  
-18'd7766,  18'd7845,  -18'd9172,  18'd3873,  -18'd550,  -18'd3240,  -18'd8040,  -18'd9208,  18'd3048,  -18'd5466,  18'd6894,  -18'd3459,  -18'd6918,  -18'd5828,  -18'd6672,  -18'd4900,  
-18'd7649,  18'd5415,  18'd4988,  18'd4292,  18'd8448,  -18'd1920,  -18'd522,  18'd4595,  -18'd3717,  -18'd5736,  -18'd9653,  -18'd7659,  18'd217,  -18'd6775,  18'd476,  18'd5675,  

18'd4867,  18'd4713,  -18'd5049,  -18'd6616,  -18'd1697,  -18'd9217,  18'd661,  18'd3521,  -18'd5012,  18'd2792,  -18'd7770,  18'd2261,  -18'd6514,  18'd5870,  -18'd8481,  -18'd5752,  
18'd6232,  18'd2420,  18'd6066,  18'd4975,  18'd6154,  -18'd4160,  -18'd2645,  -18'd11744,  -18'd2670,  -18'd8144,  -18'd11774,  18'd2689,  18'd8733,  -18'd623,  -18'd3642,  -18'd10052,  
18'd2451,  -18'd4649,  -18'd6026,  18'd1960,  18'd5045,  18'd1619,  -18'd8788,  -18'd570,  -18'd10055,  -18'd4912,  18'd7432,  18'd6300,  18'd3246,  -18'd1436,  -18'd10897,  18'd3398,  
18'd4370,  -18'd1401,  -18'd3898,  -18'd11178,  -18'd6770,  -18'd8184,  -18'd6345,  18'd4150,  -18'd6226,  18'd4830,  -18'd224,  18'd5793,  18'd3665,  -18'd3513,  18'd2351,  18'd4866,  
-18'd922,  -18'd4897,  18'd5118,  18'd5412,  -18'd6907,  -18'd10957,  18'd4986,  -18'd1438,  -18'd9320,  -18'd7488,  18'd4763,  -18'd2863,  18'd6512,  -18'd4302,  -18'd11043,  -18'd4150,  
-18'd9757,  18'd4870,  -18'd880,  18'd38,  -18'd2642,  -18'd11668,  -18'd3977,  18'd4034,  -18'd864,  -18'd2590,  18'd152,  -18'd7237,  -18'd7293,  18'd1574,  18'd2479,  -18'd4606,  
-18'd11132,  -18'd5004,  18'd33,  -18'd7553,  -18'd6253,  18'd5637,  -18'd5927,  -18'd7220,  -18'd2040,  -18'd5705,  18'd5203,  -18'd620,  -18'd8908,  -18'd8602,  -18'd6791,  -18'd8380,  
-18'd5269,  -18'd7604,  -18'd3166,  -18'd5101,  -18'd111,  18'd305,  -18'd3457,  -18'd9570,  18'd3208,  -18'd635,  -18'd2910,  -18'd2859,  -18'd1390,  -18'd3208,  -18'd12289,  -18'd5765,  
-18'd4186,  18'd5197,  -18'd5658,  18'd5272,  18'd6471,  -18'd10553,  -18'd6089,  -18'd426,  18'd5751,  -18'd3317,  -18'd9129,  -18'd1061,  -18'd4330,  18'd1993,  18'd4355,  18'd8068,  
18'd1701,  18'd1362,  -18'd248,  18'd257,  18'd2488,  -18'd4225,  -18'd1935,  18'd3947,  18'd1284,  -18'd8831,  -18'd8316,  18'd211,  -18'd4432,  18'd69,  -18'd10698,  -18'd5830,  
-18'd4776,  -18'd5039,  -18'd4198,  -18'd291,  -18'd7869,  18'd4267,  18'd5079,  -18'd6365,  -18'd8322,  -18'd3299,  18'd6093,  -18'd811,  -18'd6655,  -18'd7999,  -18'd1755,  -18'd6812,  
-18'd5601,  -18'd8901,  18'd6083,  18'd3928,  -18'd3442,  -18'd908,  18'd3959,  18'd3920,  -18'd4817,  18'd4794,  -18'd6650,  18'd5628,  -18'd5575,  -18'd6634,  -18'd9519,  18'd1094,  
18'd94,  -18'd3656,  18'd3212,  18'd3620,  18'd2489,  18'd461,  18'd3877,  -18'd10502,  -18'd8858,  18'd1395,  18'd1641,  -18'd354,  18'd6755,  -18'd1538,  -18'd262,  -18'd2516,  
18'd4117,  -18'd8204,  18'd1340,  18'd778,  18'd2694,  18'd3335,  -18'd2193,  18'd5110,  18'd1677,  18'd435,  -18'd2408,  -18'd2693,  18'd8206,  -18'd962,  -18'd11011,  -18'd8525,  
-18'd3487,  -18'd4402,  18'd2226,  18'd908,  -18'd5454,  -18'd10977,  -18'd6970,  -18'd8018,  -18'd4448,  18'd3283,  18'd406,  -18'd1804,  18'd1717,  -18'd646,  18'd5242,  -18'd8264,  
-18'd9525,  -18'd7500,  18'd1208,  18'd2705,  18'd6875,  -18'd11935,  18'd125,  18'd4626,  -18'd1475,  -18'd8265,  -18'd6615,  18'd1664,  18'd7812,  -18'd3471,  18'd253,  18'd1443,  

18'd10180,  18'd3614,  -18'd12030,  18'd6971,  -18'd6573,  -18'd23644,  -18'd17816,  18'd3346,  -18'd7048,  18'd6207,  -18'd1471,  18'd2815,  18'd7435,  -18'd8507,  -18'd16585,  -18'd1727,  
-18'd1824,  18'd25671,  -18'd1934,  18'd434,  -18'd1754,  -18'd17932,  18'd790,  18'd5587,  -18'd1487,  18'd13443,  -18'd127,  18'd6313,  18'd9842,  18'd5012,  -18'd12048,  -18'd8085,  
18'd8833,  18'd1812,  -18'd23633,  -18'd14250,  -18'd7548,  18'd6950,  18'd3502,  -18'd8087,  18'd19326,  18'd2800,  -18'd4203,  18'd17266,  -18'd3022,  -18'd4421,  18'd7227,  -18'd10361,  
18'd11648,  -18'd25765,  -18'd1160,  -18'd14310,  -18'd1607,  18'd3607,  18'd7306,  -18'd17623,  18'd3300,  -18'd22432,  18'd1434,  -18'd19995,  18'd5559,  -18'd10635,  18'd23525,  -18'd4034,  
-18'd14756,  -18'd8204,  -18'd8231,  18'd8446,  18'd3057,  -18'd4496,  -18'd6839,  -18'd3389,  18'd347,  18'd23622,  -18'd8878,  -18'd3422,  18'd9999,  18'd18280,  -18'd411,  18'd160,  
18'd3541,  18'd13019,  18'd625,  18'd14429,  18'd8394,  -18'd6108,  -18'd5547,  -18'd197,  18'd10321,  -18'd2814,  18'd679,  18'd6731,  -18'd4401,  -18'd5795,  -18'd3835,  18'd5389,  
-18'd4066,  -18'd1596,  -18'd17888,  18'd11664,  -18'd1615,  -18'd18594,  -18'd7189,  -18'd5776,  -18'd3396,  -18'd2877,  -18'd2924,  -18'd3842,  18'd9757,  18'd1705,  18'd14562,  -18'd7763,  
-18'd9373,  -18'd16734,  -18'd5732,  -18'd8048,  18'd79,  -18'd22342,  18'd18542,  18'd23358,  -18'd13437,  -18'd16964,  -18'd18176,  -18'd9754,  18'd6784,  -18'd2341,  18'd1870,  -18'd13726,  
18'd11921,  -18'd10682,  18'd1393,  -18'd16406,  -18'd891,  -18'd4232,  -18'd2777,  -18'd15317,  18'd7418,  18'd19198,  18'd8268,  18'd16471,  -18'd2646,  18'd17193,  18'd8031,  -18'd1882,  
18'd23768,  18'd11759,  -18'd6139,  18'd1465,  -18'd7123,  -18'd394,  -18'd8441,  -18'd3458,  18'd2084,  -18'd15447,  18'd13429,  18'd14584,  -18'd5911,  18'd14438,  18'd3788,  18'd4711,  
18'd2236,  -18'd5974,  18'd3603,  -18'd120,  -18'd2709,  -18'd10780,  18'd8160,  18'd7385,  -18'd12635,  18'd5082,  18'd7250,  18'd11569,  -18'd1719,  18'd5584,  -18'd6544,  -18'd4831,  
-18'd7641,  -18'd4960,  18'd1143,  18'd18048,  -18'd5294,  -18'd14028,  -18'd3705,  18'd1474,  -18'd2213,  18'd6866,  -18'd9904,  18'd10774,  18'd9587,  18'd7179,  -18'd1859,  -18'd14573,  
18'd17388,  18'd7080,  18'd11970,  18'd6321,  18'd5058,  18'd9806,  18'd11222,  18'd10480,  18'd23826,  18'd1597,  18'd2720,  18'd5928,  18'd3042,  18'd14513,  18'd13325,  -18'd9268,  
18'd15354,  18'd1523,  -18'd7662,  18'd7064,  18'd1823,  18'd7428,  18'd15697,  -18'd24845,  -18'd400,  -18'd15910,  18'd8780,  -18'd3747,  -18'd1516,  18'd11062,  -18'd780,  18'd5930,  
18'd13807,  -18'd1470,  18'd8621,  -18'd587,  -18'd1161,  18'd3234,  18'd2155,  -18'd395,  -18'd5436,  18'd14301,  -18'd5618,  18'd12444,  18'd508,  18'd1212,  -18'd7195,  18'd1437,  
18'd17169,  -18'd7719,  -18'd130,  -18'd3324,  18'd1002,  -18'd5301,  -18'd17243,  -18'd6175,  18'd16072,  18'd23448,  18'd18079,  18'd5763,  18'd6370,  18'd4929,  -18'd4231,  -18'd7843,  

-18'd39725,  18'd15550,  18'd16663,  -18'd12978,  -18'd7085,  18'd2339,  18'd12084,  18'd11061,  -18'd21686,  -18'd20393,  18'd13422,  -18'd29202,  18'd1452,  -18'd17607,  -18'd618,  18'd20565,  
-18'd20209,  18'd25590,  18'd14235,  -18'd41862,  18'd5198,  18'd17989,  18'd15267,  18'd18973,  18'd2075,  18'd1556,  -18'd3038,  -18'd13027,  -18'd5567,  -18'd1724,  18'd1409,  18'd17933,  
18'd4738,  18'd9490,  -18'd2855,  -18'd8742,  -18'd5413,  18'd16922,  -18'd11749,  -18'd7067,  18'd13833,  18'd14367,  18'd3117,  -18'd7131,  -18'd4928,  18'd5423,  18'd4633,  18'd19977,  
-18'd8119,  18'd1400,  -18'd1968,  18'd16070,  18'd4193,  18'd5519,  -18'd14710,  -18'd19301,  18'd4495,  18'd26183,  18'd24793,  18'd2961,  -18'd9435,  -18'd7512,  18'd12598,  18'd18337,  
-18'd6676,  18'd4988,  -18'd3672,  -18'd162,  -18'd6994,  18'd16318,  18'd2262,  -18'd131,  18'd19278,  -18'd2866,  -18'd3167,  -18'd10360,  18'd1067,  18'd4879,  -18'd1057,  18'd6122,  
-18'd2859,  -18'd9929,  18'd15353,  18'd926,  18'd3840,  18'd13043,  18'd6106,  -18'd6285,  18'd5348,  -18'd7273,  18'd6965,  -18'd1520,  18'd3089,  18'd5452,  -18'd11297,  18'd12154,  
18'd6626,  18'd3009,  -18'd543,  18'd10162,  18'd842,  -18'd2050,  -18'd835,  18'd9165,  18'd5550,  -18'd1345,  -18'd5684,  18'd11915,  18'd7463,  18'd5256,  18'd1383,  -18'd2696,  
-18'd1906,  18'd134,  -18'd15184,  -18'd2420,  -18'd6968,  -18'd71,  18'd15154,  18'd15754,  18'd10005,  -18'd5283,  18'd8227,  -18'd295,  -18'd544,  18'd949,  18'd11603,  -18'd6877,  
18'd14834,  -18'd17104,  18'd3548,  18'd24814,  18'd573,  18'd12122,  -18'd3990,  18'd3602,  18'd4655,  -18'd3003,  -18'd1410,  18'd909,  -18'd3754,  -18'd1783,  -18'd9591,  -18'd23712,  
18'd837,  -18'd6591,  -18'd2132,  18'd3297,  -18'd8872,  18'd1678,  18'd7244,  18'd11762,  -18'd1508,  -18'd532,  -18'd3809,  18'd3442,  18'd1638,  18'd2196,  18'd3316,  18'd8620,  
-18'd8918,  18'd9448,  18'd4391,  18'd12761,  18'd3393,  -18'd8180,  -18'd12458,  -18'd4906,  -18'd4003,  18'd7898,  18'd2991,  -18'd2984,  -18'd3336,  -18'd8525,  18'd8492,  18'd9318,  
18'd2797,  18'd1705,  -18'd6003,  18'd8619,  18'd5588,  18'd18747,  -18'd1572,  -18'd4416,  18'd7592,  -18'd6713,  18'd13791,  -18'd10794,  -18'd8258,  -18'd4001,  18'd15393,  -18'd1587,  
18'd238,  18'd668,  -18'd606,  18'd1835,  18'd1201,  -18'd2941,  -18'd5924,  18'd3297,  -18'd5006,  18'd1601,  -18'd10003,  18'd5399,  18'd632,  18'd3255,  -18'd4983,  18'd3019,  
-18'd9422,  18'd6259,  -18'd14563,  18'd6500,  -18'd4817,  -18'd9607,  -18'd14217,  18'd13751,  -18'd5323,  -18'd1305,  -18'd9280,  18'd5104,  18'd2208,  -18'd929,  18'd1821,  18'd1716,  
-18'd5651,  18'd10398,  18'd4218,  18'd7892,  18'd2610,  -18'd14809,  18'd287,  -18'd4321,  -18'd7303,  18'd6167,  18'd3109,  18'd1415,  18'd7748,  18'd3321,  -18'd6022,  18'd3045,  
18'd3521,  18'd11378,  18'd9639,  -18'd285,  -18'd8191,  -18'd783,  -18'd9106,  18'd6058,  -18'd8771,  -18'd861,  -18'd3880,  18'd4537,  18'd700,  -18'd6826,  -18'd7377,  -18'd7597,  

18'd1138,  18'd159,  -18'd70,  -18'd9731,  18'd6638,  -18'd2534,  -18'd2176,  18'd4226,  -18'd4337,  -18'd2898,  -18'd5861,  18'd436,  18'd4376,  -18'd1946,  -18'd1738,  -18'd2866,  
-18'd3186,  -18'd541,  -18'd7533,  -18'd3525,  18'd4147,  18'd2923,  18'd3302,  -18'd1287,  18'd2480,  18'd5431,  -18'd5966,  -18'd2443,  18'd8665,  18'd6363,  -18'd8795,  -18'd3396,  
-18'd9001,  -18'd407,  -18'd1527,  -18'd8967,  18'd1038,  -18'd2073,  18'd2103,  -18'd4642,  18'd1934,  18'd7864,  -18'd3903,  18'd4342,  -18'd4591,  -18'd3116,  -18'd8551,  18'd1512,  
-18'd8225,  18'd2677,  18'd801,  -18'd182,  18'd5453,  -18'd8183,  -18'd3684,  -18'd8977,  -18'd5716,  18'd3438,  -18'd5129,  18'd949,  -18'd7733,  -18'd10469,  18'd5180,  -18'd7848,  
-18'd11040,  -18'd6393,  -18'd9160,  -18'd8156,  18'd4257,  -18'd3430,  -18'd7569,  -18'd5025,  -18'd8559,  -18'd3559,  -18'd1836,  -18'd7874,  -18'd5398,  18'd6213,  18'd5670,  18'd305,  
-18'd3129,  -18'd10653,  -18'd1597,  -18'd5957,  -18'd35,  -18'd2060,  -18'd6999,  18'd2615,  -18'd10293,  -18'd7308,  -18'd8014,  -18'd999,  18'd2086,  18'd636,  -18'd8113,  -18'd8981,  
-18'd8047,  18'd4261,  -18'd6784,  18'd2583,  -18'd3262,  -18'd6422,  -18'd3919,  -18'd7871,  -18'd6767,  18'd1841,  -18'd4908,  18'd1231,  -18'd8155,  -18'd11094,  18'd1708,  -18'd4097,  
-18'd638,  -18'd4197,  18'd7345,  -18'd8156,  18'd3273,  -18'd31,  -18'd6387,  -18'd9729,  -18'd8812,  -18'd8811,  -18'd9914,  -18'd11103,  -18'd1092,  -18'd4997,  -18'd10685,  -18'd7140,  
18'd198,  18'd238,  -18'd11192,  18'd2714,  18'd3187,  -18'd52,  18'd4620,  18'd2820,  18'd2417,  -18'd2273,  -18'd6890,  -18'd9580,  -18'd6556,  -18'd11357,  -18'd41,  -18'd5795,  
-18'd3428,  -18'd2895,  18'd1444,  -18'd3703,  -18'd1936,  -18'd3531,  18'd5025,  -18'd771,  -18'd12949,  -18'd7987,  -18'd2971,  -18'd1367,  18'd7180,  18'd2589,  -18'd373,  -18'd6869,  
-18'd8117,  -18'd4705,  -18'd9303,  -18'd6350,  -18'd8200,  18'd4875,  -18'd3418,  -18'd9496,  -18'd7487,  18'd2812,  -18'd698,  18'd1952,  -18'd8091,  -18'd3187,  -18'd1205,  -18'd10472,  
-18'd9891,  18'd971,  -18'd61,  18'd1336,  -18'd7029,  18'd40,  -18'd5519,  -18'd470,  18'd374,  18'd4177,  -18'd6655,  18'd102,  18'd1698,  -18'd8075,  -18'd1548,  -18'd350,  
-18'd8204,  -18'd9096,  18'd512,  -18'd3145,  -18'd6912,  -18'd9145,  -18'd10216,  -18'd10,  18'd3977,  -18'd11784,  18'd6269,  -18'd3776,  -18'd6471,  18'd1607,  -18'd3940,  -18'd7708,  
18'd5251,  -18'd1980,  -18'd6549,  18'd2446,  18'd7751,  -18'd6218,  18'd3242,  -18'd5695,  -18'd7870,  -18'd8318,  -18'd6933,  -18'd10757,  18'd858,  18'd6780,  -18'd2392,  18'd100,  
-18'd1518,  -18'd3552,  18'd3074,  18'd2821,  18'd5923,  -18'd7722,  -18'd6940,  18'd4364,  18'd3918,  -18'd6373,  18'd4485,  -18'd5854,  18'd1340,  -18'd10946,  -18'd2300,  -18'd9224,  
18'd967,  -18'd10354,  18'd384,  18'd886,  -18'd8265,  -18'd11545,  18'd1528,  18'd3944,  18'd3602,  18'd5410,  -18'd7045,  -18'd7660,  -18'd5567,  18'd5326,  -18'd4048,  18'd1592,  

-18'd6442,  -18'd531,  18'd334,  -18'd2319,  -18'd6537,  -18'd4467,  18'd10798,  18'd3984,  18'd6046,  18'd17854,  18'd4535,  -18'd5094,  18'd1211,  -18'd5427,  18'd21546,  -18'd13417,  
18'd17999,  -18'd3574,  18'd5139,  18'd18794,  18'd734,  18'd98,  18'd8270,  18'd11606,  18'd13261,  18'd10546,  18'd14431,  -18'd6297,  -18'd11134,  -18'd18459,  18'd24586,  18'd2372,  
18'd12507,  18'd4999,  18'd10779,  -18'd5040,  -18'd2710,  18'd10529,  18'd14876,  18'd13106,  -18'd1858,  -18'd21044,  18'd11551,  -18'd6284,  -18'd11538,  -18'd19430,  18'd12599,  -18'd6320,  
-18'd18546,  18'd15107,  18'd21310,  18'd15807,  -18'd6277,  -18'd9339,  -18'd13883,  18'd17252,  -18'd4579,  -18'd1203,  -18'd19787,  -18'd13490,  -18'd12365,  -18'd4890,  18'd1206,  -18'd2281,  
18'd1475,  18'd5196,  18'd8365,  -18'd18619,  -18'd2219,  -18'd1628,  18'd3371,  18'd13420,  18'd13691,  18'd7043,  18'd10611,  18'd3189,  -18'd7103,  -18'd4048,  18'd10363,  18'd3,  
-18'd3555,  18'd13621,  18'd5078,  -18'd5917,  -18'd6192,  -18'd4781,  18'd22538,  18'd10501,  -18'd5913,  18'd10469,  -18'd4528,  18'd5804,  -18'd1588,  18'd8236,  18'd2029,  -18'd6880,  
18'd3868,  18'd4022,  18'd22479,  -18'd3213,  -18'd1166,  18'd17861,  18'd15601,  18'd10865,  18'd4743,  -18'd18423,  -18'd4609,  18'd4468,  18'd3772,  -18'd5380,  -18'd8795,  18'd19709,  
-18'd16268,  18'd9859,  18'd12986,  18'd16011,  18'd7605,  -18'd3520,  -18'd13819,  18'd1653,  -18'd5866,  -18'd6286,  -18'd12946,  -18'd1023,  -18'd4647,  18'd6469,  18'd1566,  18'd38494,  
18'd14638,  -18'd2828,  -18'd2442,  18'd8225,  18'd8698,  18'd4484,  -18'd871,  18'd15529,  -18'd5850,  18'd16402,  -18'd3813,  18'd13681,  -18'd10317,  18'd3469,  -18'd6536,  -18'd5207,  
18'd2254,  18'd281,  -18'd11003,  18'd11569,  18'd1795,  18'd4128,  -18'd2214,  18'd8266,  -18'd4067,  18'd14154,  18'd8134,  18'd25024,  -18'd11870,  18'd4463,  18'd1399,  18'd13066,  
18'd2558,  -18'd6000,  18'd22207,  18'd11015,  -18'd3715,  18'd10104,  -18'd18515,  18'd4087,  18'd6674,  18'd9545,  18'd6557,  18'd16641,  18'd2927,  18'd6519,  -18'd9920,  -18'd3236,  
18'd485,  18'd7623,  -18'd9700,  18'd10444,  -18'd5289,  18'd5248,  18'd3245,  -18'd10373,  -18'd4500,  -18'd17985,  -18'd19598,  -18'd9806,  -18'd9880,  18'd283,  18'd5473,  -18'd3358,  
-18'd3253,  -18'd10165,  -18'd20487,  -18'd8468,  18'd4156,  -18'd8822,  -18'd8632,  -18'd4608,  -18'd4733,  18'd17458,  -18'd9755,  18'd1149,  -18'd3170,  18'd12830,  18'd9716,  -18'd8315,  
18'd9770,  18'd9414,  -18'd3355,  -18'd2201,  18'd5800,  -18'd7531,  -18'd14505,  -18'd4540,  -18'd6751,  18'd23132,  -18'd4142,  -18'd528,  18'd1537,  18'd11007,  -18'd4477,  -18'd806,  
-18'd4197,  18'd16904,  -18'd9079,  -18'd4120,  18'd8373,  18'd6739,  -18'd15323,  -18'd9170,  -18'd1309,  -18'd2466,  18'd729,  18'd5863,  -18'd7973,  18'd9581,  -18'd10451,  -18'd6378,  
18'd6444,  -18'd1900,  -18'd20190,  18'd9493,  -18'd9048,  18'd11577,  -18'd4447,  18'd6079,  18'd3418,  -18'd1115,  18'd12069,  18'd760,  18'd3702,  18'd3744,  -18'd2726,  -18'd13691,  

18'd33347,  18'd2399,  -18'd1898,  18'd24407,  -18'd1062,  18'd8213,  -18'd4980,  -18'd8232,  18'd17087,  18'd6281,  18'd4190,  18'd17984,  -18'd10171,  18'd16434,  -18'd9353,  18'd19676,  
-18'd13,  18'd3732,  18'd5870,  18'd17252,  -18'd2688,  -18'd5641,  -18'd1259,  -18'd10282,  18'd1231,  -18'd35947,  -18'd1381,  -18'd1304,  -18'd12858,  -18'd9982,  -18'd2566,  18'd22765,  
-18'd10529,  18'd4404,  18'd4273,  18'd2818,  -18'd2834,  -18'd3363,  18'd16814,  -18'd5269,  -18'd11371,  -18'd40389,  18'd11985,  -18'd23002,  -18'd12805,  -18'd18288,  -18'd13568,  18'd8439,  
-18'd311,  -18'd17784,  18'd18393,  -18'd11592,  -18'd8170,  -18'd7592,  18'd24341,  -18'd4474,  -18'd18475,  -18'd12595,  -18'd22755,  -18'd45379,  -18'd4229,  -18'd15972,  -18'd16794,  -18'd1328,  
18'd18701,  18'd3464,  -18'd4045,  18'd29306,  18'd8032,  18'd4869,  -18'd3710,  -18'd8825,  18'd3145,  18'd9750,  18'd9008,  18'd15061,  -18'd5491,  18'd4411,  18'd5158,  18'd1364,  
-18'd19775,  18'd16446,  -18'd690,  18'd21535,  18'd5809,  18'd4501,  -18'd14655,  -18'd1415,  18'd5969,  -18'd9981,  -18'd3347,  18'd1822,  -18'd1471,  -18'd3393,  -18'd179,  -18'd4533,  
-18'd7033,  18'd3633,  18'd9124,  -18'd6728,  18'd7110,  18'd4439,  18'd8044,  -18'd931,  18'd22938,  -18'd4913,  18'd8244,  18'd3780,  -18'd580,  18'd9400,  -18'd23134,  18'd19397,  
18'd4874,  -18'd8619,  18'd9345,  18'd3916,  -18'd3391,  18'd10907,  18'd3697,  -18'd3065,  18'd6121,  18'd849,  -18'd668,  -18'd6941,  18'd4004,  18'd9818,  -18'd4309,  18'd11838,  
-18'd9985,  18'd14989,  18'd4058,  -18'd3514,  -18'd5135,  -18'd5113,  -18'd15176,  18'd12770,  18'd1304,  18'd7741,  -18'd1406,  18'd10828,  -18'd3423,  18'd8359,  18'd10689,  18'd18549,  
-18'd14099,  18'd14324,  -18'd8492,  -18'd8689,  -18'd437,  -18'd2118,  -18'd7458,  18'd10874,  -18'd4744,  18'd231,  18'd7273,  18'd528,  -18'd6003,  18'd8697,  -18'd2559,  18'd7278,  
-18'd11409,  18'd11014,  18'd1965,  -18'd3021,  18'd6868,  -18'd1154,  18'd9980,  18'd3967,  18'd5064,  18'd1554,  -18'd8230,  -18'd2272,  -18'd889,  18'd7213,  -18'd12861,  18'd15436,  
18'd10769,  18'd5990,  18'd274,  18'd1035,  18'd4547,  -18'd4665,  -18'd1917,  18'd7468,  -18'd10648,  18'd25088,  -18'd3572,  18'd5789,  -18'd12744,  18'd5896,  -18'd951,  18'd5711,  
18'd6180,  -18'd12875,  18'd707,  -18'd11224,  18'd2266,  -18'd15175,  18'd1290,  -18'd1245,  18'd631,  18'd11454,  18'd7079,  18'd2394,  -18'd1516,  -18'd72,  18'd12278,  -18'd12089,  
18'd3489,  -18'd8168,  -18'd9487,  -18'd8696,  -18'd2612,  -18'd5923,  -18'd10303,  18'd2263,  -18'd4992,  18'd5676,  18'd11800,  -18'd1849,  -18'd307,  18'd9109,  -18'd1682,  -18'd11772,  
18'd3434,  -18'd18460,  -18'd6653,  18'd5546,  18'd8436,  18'd1533,  18'd7858,  18'd1099,  -18'd2606,  18'd13931,  -18'd567,  -18'd787,  18'd2546,  -18'd14358,  18'd11987,  -18'd14117,  
-18'd8309,  18'd955,  -18'd3714,  18'd18019,  -18'd3481,  18'd4893,  18'd13818,  18'd3085,  -18'd10661,  18'd19830,  18'd15274,  18'd4553,  18'd1752,  18'd12649,  18'd6923,  18'd11675,  

-18'd5917,  18'd3766,  -18'd8227,  -18'd3596,  18'd2365,  -18'd9810,  -18'd886,  -18'd8865,  -18'd6257,  -18'd282,  18'd4580,  -18'd978,  18'd5045,  -18'd8084,  -18'd8169,  -18'd1553,  
-18'd3104,  -18'd10184,  -18'd7275,  18'd984,  18'd2136,  -18'd1665,  -18'd6260,  -18'd584,  -18'd3233,  18'd4870,  18'd3382,  -18'd10097,  18'd160,  18'd6361,  -18'd5616,  18'd6928,  
-18'd4243,  18'd4346,  18'd5740,  -18'd2684,  -18'd5623,  18'd8901,  -18'd7675,  -18'd368,  18'd2094,  -18'd4317,  -18'd10431,  -18'd1245,  18'd3337,  18'd5127,  18'd998,  -18'd2630,  
-18'd6860,  -18'd1842,  -18'd6034,  -18'd5025,  18'd4461,  -18'd5480,  -18'd4529,  18'd230,  18'd947,  -18'd3131,  18'd1593,  -18'd4907,  -18'd3124,  -18'd4997,  -18'd2238,  -18'd9660,  
18'd2622,  -18'd5962,  18'd679,  18'd2712,  18'd4213,  -18'd1770,  18'd3332,  -18'd2223,  18'd6306,  18'd7385,  18'd564,  18'd6510,  -18'd1890,  -18'd6150,  18'd5458,  -18'd5242,  
18'd2905,  18'd5290,  18'd1585,  -18'd3651,  18'd4212,  18'd1792,  18'd2571,  -18'd9116,  -18'd8530,  18'd1050,  18'd5977,  18'd2145,  18'd153,  -18'd6921,  18'd2695,  18'd5537,  
18'd330,  18'd111,  18'd3720,  -18'd6553,  -18'd5970,  -18'd141,  -18'd2179,  -18'd4550,  -18'd9981,  -18'd13050,  -18'd1829,  -18'd6726,  -18'd658,  -18'd11106,  18'd4474,  18'd6984,  
-18'd5110,  -18'd457,  18'd101,  18'd1976,  18'd956,  18'd2653,  18'd1951,  18'd1710,  -18'd2872,  18'd1174,  18'd1688,  -18'd10772,  -18'd1459,  -18'd9948,  -18'd11358,  18'd2995,  
-18'd6226,  -18'd5577,  -18'd4413,  -18'd4891,  18'd6124,  18'd3000,  18'd429,  -18'd2805,  -18'd340,  18'd6445,  -18'd6150,  -18'd9971,  -18'd4809,  18'd371,  -18'd429,  -18'd4729,  
-18'd6114,  18'd254,  -18'd10866,  -18'd8578,  -18'd861,  18'd3461,  18'd4418,  -18'd8157,  -18'd2360,  18'd535,  18'd2954,  -18'd6063,  18'd3407,  18'd849,  18'd3202,  -18'd7376,  
18'd728,  18'd8258,  -18'd634,  -18'd1411,  -18'd6738,  -18'd8852,  -18'd4996,  -18'd9468,  18'd6387,  -18'd10961,  -18'd2173,  -18'd7725,  18'd1148,  -18'd6243,  -18'd11756,  18'd802,  
18'd4248,  18'd1326,  -18'd10485,  18'd2394,  18'd5598,  -18'd6942,  -18'd4353,  -18'd1374,  -18'd7080,  18'd2188,  -18'd11017,  -18'd2296,  -18'd7279,  18'd228,  18'd3215,  18'd6643,  
18'd1234,  -18'd5371,  -18'd11066,  18'd4278,  18'd4539,  18'd561,  -18'd857,  -18'd5692,  -18'd7669,  -18'd3627,  -18'd619,  -18'd1023,  -18'd1588,  18'd3728,  18'd2727,  18'd7822,  
-18'd4898,  -18'd2433,  -18'd6653,  18'd1222,  -18'd4387,  -18'd10829,  -18'd880,  18'd2243,  -18'd8441,  18'd5207,  -18'd3773,  -18'd8359,  18'd7603,  18'd3008,  -18'd6311,  18'd4524,  
18'd3755,  -18'd408,  18'd7247,  -18'd3006,  18'd2578,  -18'd8237,  -18'd9773,  18'd7212,  18'd1004,  -18'd4621,  -18'd9579,  -18'd1716,  18'd2876,  18'd1420,  -18'd5474,  -18'd6362,  
18'd6360,  -18'd12360,  -18'd11723,  -18'd3352,  18'd117,  -18'd11066,  -18'd8091,  18'd3098,  18'd860,  -18'd9104,  -18'd11380,  -18'd58,  -18'd2818,  18'd3152,  -18'd4552,  -18'd2795,  

-18'd11280,  -18'd30073,  18'd1651,  18'd13031,  18'd4292,  -18'd2752,  18'd12151,  -18'd2394,  -18'd9203,  18'd20857,  18'd9465,  -18'd11975,  18'd8141,  -18'd24576,  18'd16905,  -18'd24263,  
18'd14624,  18'd8298,  18'd8979,  -18'd2821,  18'd3504,  18'd3288,  18'd31305,  18'd11282,  18'd22732,  18'd14890,  18'd14801,  -18'd3007,  18'd7601,  -18'd20703,  18'd22507,  -18'd13757,  
18'd3971,  18'd2056,  18'd833,  -18'd12898,  -18'd5083,  18'd2536,  18'd3233,  18'd5995,  18'd21004,  -18'd16113,  -18'd13046,  18'd6244,  18'd6301,  -18'd987,  18'd3177,  -18'd3504,  
18'd8947,  -18'd3549,  18'd9897,  -18'd10614,  18'd4387,  18'd4855,  18'd21538,  18'd4887,  18'd746,  -18'd20951,  -18'd2159,  -18'd2204,  -18'd6296,  -18'd14881,  18'd1533,  -18'd15120,  
-18'd12384,  18'd688,  18'd8228,  18'd4973,  -18'd4817,  -18'd8632,  18'd8476,  18'd19756,  -18'd1050,  -18'd4862,  18'd1350,  18'd1288,  18'd4786,  18'd2390,  -18'd3717,  -18'd13802,  
18'd4020,  18'd22298,  18'd21475,  -18'd19211,  -18'd2865,  18'd3538,  -18'd9583,  18'd23047,  -18'd1481,  -18'd9406,  18'd12438,  18'd15668,  -18'd3079,  18'd6976,  18'd8327,  18'd3665,  
18'd2332,  18'd19692,  -18'd2738,  -18'd19,  18'd5352,  18'd9246,  -18'd20458,  18'd5085,  18'd362,  -18'd11262,  -18'd7564,  18'd594,  -18'd5714,  18'd20409,  18'd6734,  18'd5066,  
-18'd240,  18'd28656,  18'd3493,  18'd6986,  18'd4636,  -18'd8679,  -18'd5990,  18'd16970,  -18'd18918,  -18'd5052,  -18'd29416,  18'd10599,  18'd6759,  18'd2790,  -18'd1950,  18'd8558,  
-18'd1496,  18'd8514,  18'd6223,  -18'd14303,  18'd809,  -18'd5142,  -18'd6365,  18'd21,  -18'd3970,  18'd10838,  18'd3819,  18'd6228,  18'd9325,  18'd2733,  -18'd4061,  -18'd10525,  
18'd548,  18'd20092,  -18'd10378,  -18'd10007,  18'd108,  -18'd5265,  -18'd19635,  18'd21177,  18'd3755,  -18'd1203,  -18'd7109,  18'd8545,  18'd8642,  18'd24035,  -18'd9145,  18'd10522,  
-18'd7531,  18'd14317,  -18'd2145,  18'd6316,  -18'd5835,  -18'd11561,  18'd501,  18'd5234,  -18'd6824,  18'd12048,  18'd10439,  18'd2183,  -18'd1700,  18'd16744,  -18'd3214,  18'd25,  
18'd9014,  18'd18242,  -18'd6905,  18'd25743,  18'd6108,  -18'd8456,  -18'd5520,  -18'd11406,  18'd12446,  18'd5916,  -18'd1395,  18'd3448,  18'd6489,  18'd12063,  -18'd6082,  18'd26126,  
18'd7377,  18'd1048,  -18'd11944,  -18'd4930,  -18'd7398,  -18'd13304,  -18'd7259,  18'd7725,  -18'd3734,  18'd16432,  18'd996,  18'd6568,  18'd4096,  18'd6104,  -18'd1791,  18'd8325,  
18'd9163,  18'd7542,  -18'd9689,  18'd2974,  18'd7595,  -18'd17772,  -18'd5324,  -18'd15846,  -18'd12405,  -18'd2125,  18'd457,  -18'd12959,  18'd6418,  18'd9819,  -18'd4378,  18'd3758,  
18'd9929,  -18'd3478,  18'd2213,  18'd240,  18'd4954,  18'd13157,  18'd4469,  -18'd15047,  -18'd10315,  18'd4326,  18'd2899,  18'd14895,  -18'd7659,  18'd10505,  18'd6101,  -18'd14966,  
18'd4848,  -18'd20541,  -18'd2516,  18'd6939,  18'd2365,  18'd10626,  -18'd3845,  -18'd14025,  18'd21195,  -18'd7689,  18'd4124,  -18'd5460,  18'd5780,  18'd1007,  18'd2822,  -18'd7910,  

-18'd24554,  18'd22029,  -18'd11805,  18'd10154,  18'd8151,  -18'd18919,  -18'd1513,  18'd9381,  -18'd21059,  18'd193,  18'd1830,  -18'd14191,  -18'd7822,  -18'd30230,  -18'd691,  -18'd11488,  
-18'd8958,  -18'd2084,  -18'd4759,  -18'd15050,  -18'd1535,  18'd744,  18'd7650,  18'd1887,  -18'd11346,  -18'd8840,  -18'd278,  -18'd15226,  18'd3078,  -18'd14643,  18'd10706,  -18'd6825,  
18'd4634,  -18'd11273,  -18'd1959,  -18'd22670,  -18'd6177,  18'd12652,  18'd15960,  -18'd7563,  18'd3345,  18'd4174,  -18'd4347,  -18'd7769,  -18'd10227,  -18'd9612,  18'd12599,  -18'd8570,  
18'd13486,  -18'd1762,  18'd13725,  -18'd10089,  18'd5589,  18'd1193,  18'd294,  -18'd8317,  18'd9725,  -18'd24,  18'd4503,  -18'd13268,  -18'd695,  -18'd8882,  -18'd903,  -18'd3600,  
-18'd15374,  18'd16060,  -18'd1389,  18'd11772,  -18'd4409,  18'd1465,  18'd1084,  18'd9178,  18'd1610,  18'd15044,  -18'd4636,  18'd6326,  -18'd756,  -18'd31,  -18'd2970,  18'd10253,  
-18'd7558,  18'd13832,  18'd2394,  -18'd1827,  -18'd2684,  18'd2238,  -18'd7048,  18'd20447,  -18'd12816,  -18'd6879,  18'd3640,  -18'd1595,  18'd5239,  -18'd7942,  18'd5362,  18'd14010,  
18'd6922,  18'd36111,  18'd17903,  -18'd6814,  18'd564,  18'd10720,  18'd15786,  18'd27953,  18'd4084,  -18'd8663,  18'd6379,  -18'd13711,  -18'd7561,  18'd2260,  18'd12479,  18'd2110,  
18'd6029,  18'd6699,  18'd8823,  18'd7693,  18'd3602,  18'd23036,  18'd10592,  18'd22014,  18'd10803,  18'd1349,  -18'd196,  18'd1143,  18'd508,  18'd5583,  -18'd10710,  18'd2431,  
-18'd16433,  18'd4389,  18'd4886,  18'd7254,  -18'd7684,  18'd10274,  -18'd3011,  -18'd7011,  18'd2160,  18'd17103,  18'd28,  18'd8707,  -18'd11168,  18'd19141,  -18'd16205,  18'd23931,  
-18'd4116,  18'd12394,  -18'd6225,  18'd38798,  18'd2938,  18'd3054,  -18'd1486,  -18'd4348,  18'd9628,  18'd2935,  18'd10647,  -18'd5253,  -18'd10427,  18'd15213,  -18'd9457,  18'd16774,  
-18'd1388,  18'd28931,  18'd12055,  18'd12910,  18'd1512,  -18'd5655,  18'd14889,  18'd13589,  18'd2026,  18'd5024,  18'd10670,  -18'd3918,  18'd174,  18'd2953,  -18'd6178,  18'd10705,  
18'd6504,  18'd3861,  18'd14273,  18'd937,  -18'd5603,  18'd10192,  18'd10747,  -18'd3583,  18'd7342,  18'd20653,  18'd4454,  -18'd5272,  -18'd5207,  18'd12083,  -18'd4296,  18'd7138,  
-18'd7428,  -18'd8734,  18'd2159,  18'd14488,  -18'd3825,  -18'd1582,  -18'd13129,  -18'd13199,  18'd5977,  18'd6119,  -18'd8225,  18'd17667,  18'd4588,  18'd10345,  18'd972,  -18'd1925,  
18'd14032,  18'd5532,  -18'd9429,  18'd30168,  -18'd2179,  18'd5756,  18'd3033,  -18'd26223,  18'd5387,  -18'd11666,  -18'd1050,  -18'd8391,  -18'd3531,  18'd15376,  18'd4224,  -18'd2000,  
-18'd1512,  18'd9504,  -18'd7025,  18'd13430,  18'd4067,  -18'd9646,  -18'd7716,  -18'd13065,  -18'd309,  -18'd12212,  18'd5435,  -18'd7771,  18'd1838,  -18'd1163,  18'd5537,  18'd5257,  
-18'd6802,  18'd4194,  18'd4967,  -18'd5588,  18'd4287,  18'd23186,  18'd5765,  18'd5338,  18'd9244,  -18'd5888,  18'd10031,  18'd6000,  -18'd2335,  18'd13921,  -18'd13655,  18'd5497,  

18'd17765,  -18'd4514,  -18'd3129,  18'd9859,  -18'd7926,  -18'd9777,  -18'd5843,  -18'd910,  18'd4216,  18'd13960,  18'd2008,  18'd11857,  -18'd8484,  18'd4014,  18'd15790,  -18'd6836,  
-18'd10203,  18'd8216,  18'd7924,  -18'd1800,  18'd3876,  18'd16632,  18'd2948,  18'd7124,  18'd16906,  -18'd81,  18'd2911,  18'd17250,  18'd4919,  -18'd9839,  18'd1003,  -18'd8912,  
-18'd5135,  18'd12994,  18'd6748,  -18'd6391,  18'd3221,  18'd10581,  18'd15037,  -18'd7853,  -18'd3801,  -18'd29715,  18'd14209,  -18'd10121,  -18'd9607,  18'd6339,  -18'd10606,  18'd8553,  
-18'd7811,  18'd16581,  18'd4146,  18'd7496,  -18'd7429,  -18'd6031,  -18'd1487,  18'd7318,  18'd5701,  -18'd2352,  -18'd22709,  -18'd23905,  -18'd4631,  18'd5585,  -18'd17088,  18'd6313,  
-18'd469,  18'd17645,  18'd8410,  18'd8499,  18'd5835,  -18'd11711,  -18'd2344,  18'd16303,  -18'd5213,  -18'd7259,  -18'd368,  -18'd8160,  -18'd1589,  -18'd6614,  18'd9556,  18'd18803,  
-18'd11054,  18'd12088,  -18'd774,  -18'd3933,  -18'd4566,  18'd8522,  18'd10802,  18'd5873,  -18'd3023,  -18'd4064,  18'd953,  -18'd8120,  -18'd9750,  18'd3038,  -18'd6053,  -18'd7222,  
-18'd3310,  -18'd5120,  18'd18675,  -18'd8661,  18'd4656,  18'd9734,  18'd1321,  -18'd704,  18'd9166,  -18'd4330,  -18'd3196,  -18'd14963,  -18'd6952,  18'd5194,  -18'd20720,  18'd12010,  
18'd7263,  -18'd9934,  -18'd10032,  18'd10014,  18'd5720,  18'd7618,  -18'd4175,  -18'd16468,  18'd8680,  18'd9069,  -18'd5436,  18'd2929,  18'd4578,  18'd16374,  -18'd7440,  18'd16970,  
18'd5583,  -18'd951,  18'd9913,  18'd16244,  18'd4666,  -18'd19608,  18'd5428,  18'd16118,  18'd2062,  18'd3961,  18'd4815,  18'd6887,  18'd1088,  18'd4118,  18'd5117,  18'd7983,  
-18'd6490,  18'd14875,  -18'd8624,  -18'd23593,  -18'd3359,  -18'd528,  -18'd3172,  18'd6447,  18'd4523,  -18'd3317,  18'd9908,  18'd11510,  18'd6344,  18'd13853,  -18'd11389,  -18'd5,  
-18'd8303,  18'd3574,  18'd2608,  18'd2089,  -18'd2987,  -18'd2037,  18'd9980,  18'd11679,  18'd8320,  -18'd1642,  18'd751,  -18'd6042,  18'd549,  -18'd5514,  18'd606,  18'd3993,  
18'd15929,  18'd172,  -18'd2530,  18'd1009,  -18'd3026,  18'd4764,  18'd11626,  18'd3521,  -18'd183,  -18'd9770,  -18'd356,  18'd1129,  -18'd3351,  -18'd1093,  18'd4411,  -18'd9569,  
-18'd243,  -18'd12605,  -18'd10194,  18'd11080,  -18'd8611,  -18'd6252,  18'd9838,  18'd3153,  18'd777,  18'd16191,  18'd1356,  -18'd4851,  -18'd1009,  -18'd15418,  18'd14885,  -18'd4951,  
18'd17209,  -18'd9663,  18'd5230,  -18'd27837,  -18'd8646,  18'd190,  -18'd2106,  18'd5868,  18'd1941,  18'd5840,  18'd8378,  18'd8605,  -18'd9759,  -18'd8000,  18'd7,  -18'd7392,  
-18'd6034,  -18'd9526,  18'd6275,  18'd8039,  -18'd8233,  -18'd4511,  -18'd4283,  18'd14298,  18'd2365,  -18'd192,  -18'd1150,  -18'd3695,  18'd2189,  18'd4806,  18'd7433,  18'd6413,  
-18'd212,  -18'd4614,  -18'd1103,  18'd5739,  -18'd6613,  -18'd4593,  18'd11103,  18'd11367,  18'd582,  18'd2426,  18'd14073,  18'd9215,  -18'd5987,  18'd214,  -18'd3178,  18'd1702,  

-18'd4718,  18'd15824,  18'd6762,  18'd8310,  18'd3225,  -18'd12808,  -18'd3278,  18'd2380,  -18'd8717,  -18'd1723,  -18'd7203,  -18'd7705,  18'd10139,  18'd10486,  18'd2747,  18'd8873,  
-18'd7557,  18'd538,  18'd2104,  18'd10615,  18'd4542,  -18'd890,  -18'd11287,  18'd5684,  -18'd1718,  18'd20665,  18'd8779,  18'd6369,  18'd689,  18'd4357,  18'd784,  -18'd9449,  
18'd8192,  -18'd1751,  -18'd849,  18'd9375,  -18'd3075,  18'd15963,  -18'd1840,  -18'd91,  18'd13639,  -18'd4765,  18'd7068,  18'd11317,  -18'd4373,  18'd7908,  -18'd5421,  -18'd4854,  
18'd4211,  -18'd12943,  -18'd8172,  18'd3777,  18'd7743,  -18'd1760,  18'd12481,  18'd14075,  18'd15728,  -18'd8943,  -18'd27300,  -18'd9431,  18'd3086,  -18'd9071,  18'd6655,  -18'd2444,  
-18'd8023,  -18'd1768,  -18'd541,  -18'd7325,  -18'd5211,  -18'd1587,  -18'd1360,  -18'd6732,  -18'd1702,  -18'd11036,  18'd5426,  18'd1195,  18'd1970,  -18'd2185,  -18'd707,  18'd11130,  
18'd9331,  -18'd15108,  18'd4379,  18'd5525,  18'd1954,  -18'd12758,  18'd6343,  -18'd18447,  -18'd928,  18'd579,  18'd5213,  -18'd5367,  -18'd2986,  -18'd6676,  18'd7238,  18'd3948,  
-18'd9865,  -18'd15675,  -18'd652,  18'd9357,  18'd5915,  18'd555,  18'd698,  -18'd9468,  -18'd2988,  -18'd2772,  -18'd11430,  -18'd14809,  18'd1077,  18'd6910,  18'd9177,  18'd263,  
-18'd11120,  18'd5657,  -18'd21376,  18'd21053,  18'd59,  -18'd11560,  -18'd1942,  18'd3206,  -18'd3213,  -18'd11003,  -18'd16586,  -18'd14137,  18'd3879,  -18'd5827,  18'd3184,  -18'd9893,  
18'd17627,  18'd1668,  18'd5462,  18'd10869,  -18'd7500,  18'd4338,  -18'd3710,  -18'd2030,  18'd1172,  18'd2648,  -18'd2919,  18'd7418,  18'd12163,  18'd1891,  -18'd2527,  -18'd13342,  
-18'd7124,  -18'd2866,  18'd5711,  18'd901,  -18'd794,  18'd406,  18'd12692,  -18'd9339,  18'd4500,  18'd1698,  18'd9651,  -18'd6895,  18'd1220,  18'd3414,  -18'd9973,  18'd11048,  
18'd4588,  -18'd8650,  -18'd2303,  18'd1434,  18'd6363,  -18'd6751,  18'd15814,  -18'd9471,  -18'd6550,  -18'd5421,  -18'd5766,  18'd5377,  18'd3945,  18'd13144,  -18'd6586,  18'd2167,  
18'd1942,  18'd6760,  -18'd20584,  18'd22369,  -18'd4082,  18'd3474,  18'd15856,  -18'd18845,  18'd3455,  -18'd12241,  -18'd25922,  18'd1875,  18'd12126,  -18'd4896,  18'd2724,  -18'd1414,  
18'd2556,  18'd15008,  -18'd1068,  18'd34897,  -18'd2320,  18'd7333,  18'd4572,  18'd19428,  -18'd14866,  18'd15613,  -18'd5941,  18'd13777,  -18'd76,  18'd7743,  -18'd12521,  -18'd4001,  
-18'd4719,  -18'd5026,  18'd12000,  -18'd9114,  18'd1619,  18'd8440,  18'd12107,  18'd11176,  -18'd3173,  18'd1005,  18'd12024,  18'd2932,  18'd8584,  -18'd4839,  -18'd1590,  -18'd617,  
18'd13890,  -18'd6491,  18'd6309,  -18'd5611,  -18'd5775,  18'd7422,  18'd18000,  -18'd20646,  18'd57,  -18'd10048,  -18'd7738,  18'd12270,  18'd3319,  -18'd1595,  -18'd2161,  -18'd40,  
18'd12132,  -18'd24616,  18'd4798,  18'd3424,  18'd2270,  18'd26666,  18'd3527,  -18'd23825,  18'd23737,  18'd4585,  -18'd1952,  18'd4658,  18'd1907,  -18'd1200,  -18'd1090,  -18'd10465,  

-18'd1185,  -18'd3611,  18'd1806,  -18'd8365,  -18'd871,  18'd244,  18'd5995,  18'd3068,  -18'd2413,  18'd2803,  -18'd6568,  -18'd1065,  -18'd1249,  -18'd4640,  -18'd11022,  -18'd8031,  
18'd2140,  18'd1296,  18'd44,  18'd108,  -18'd2033,  18'd1876,  -18'd12650,  18'd3766,  18'd7383,  -18'd1133,  18'd1126,  -18'd240,  -18'd7230,  -18'd2575,  -18'd4317,  -18'd3442,  
18'd6220,  -18'd3424,  -18'd2984,  18'd2217,  -18'd8444,  18'd3666,  -18'd10797,  18'd4410,  -18'd6908,  18'd3270,  18'd1366,  18'd428,  18'd3003,  18'd6809,  18'd1991,  18'd5361,  
-18'd8884,  -18'd8282,  -18'd7861,  18'd589,  18'd6433,  -18'd10855,  -18'd355,  -18'd181,  -18'd11272,  -18'd11145,  18'd696,  18'd662,  -18'd1119,  -18'd6013,  18'd5156,  -18'd10871,  
18'd7394,  -18'd858,  18'd6188,  -18'd7410,  18'd5546,  -18'd899,  18'd249,  18'd2351,  -18'd7539,  18'd5430,  -18'd98,  18'd8247,  -18'd4547,  -18'd9245,  18'd4122,  -18'd2609,  
18'd3798,  18'd3535,  -18'd2713,  -18'd5471,  18'd2821,  -18'd9683,  18'd2474,  18'd1951,  -18'd2924,  -18'd8833,  18'd894,  -18'd489,  18'd1509,  -18'd5017,  18'd3932,  -18'd11568,  
-18'd6301,  -18'd8204,  18'd1099,  -18'd3190,  -18'd3137,  -18'd2932,  18'd1968,  -18'd154,  -18'd6166,  -18'd14399,  -18'd10520,  -18'd6094,  18'd7139,  -18'd4368,  -18'd4183,  -18'd13754,  
-18'd5742,  18'd9187,  18'd8416,  -18'd11956,  18'd2528,  -18'd682,  -18'd6109,  -18'd4126,  18'd3466,  18'd770,  18'd5212,  18'd2717,  -18'd8062,  18'd145,  -18'd6276,  18'd1678,  
18'd8260,  -18'd2031,  -18'd1619,  -18'd9032,  -18'd3302,  18'd322,  -18'd2377,  -18'd9231,  18'd6578,  -18'd9773,  -18'd6886,  18'd3548,  18'd5121,  -18'd130,  -18'd8646,  18'd7967,  
18'd4789,  -18'd2774,  -18'd6864,  -18'd4829,  -18'd8108,  -18'd1056,  -18'd2601,  -18'd3288,  -18'd7526,  -18'd117,  18'd3890,  -18'd773,  18'd4285,  -18'd8117,  -18'd10143,  -18'd7741,  
18'd3798,  -18'd7342,  -18'd7278,  18'd1351,  -18'd3193,  -18'd9412,  -18'd7898,  18'd7269,  -18'd8144,  -18'd9440,  -18'd5405,  -18'd8224,  -18'd1335,  -18'd12425,  -18'd11925,  -18'd8069,  
-18'd8050,  -18'd1190,  18'd2193,  -18'd4752,  18'd6012,  -18'd3182,  -18'd11049,  18'd8541,  -18'd6662,  18'd807,  18'd4000,  -18'd7632,  18'd5677,  -18'd6617,  -18'd15073,  18'd4820,  
18'd104,  -18'd2127,  -18'd6308,  18'd2469,  18'd7853,  -18'd3416,  18'd173,  18'd4476,  -18'd7343,  -18'd8098,  18'd10,  18'd3417,  18'd8828,  18'd9010,  -18'd9123,  -18'd2294,  
-18'd4317,  18'd7488,  18'd6414,  -18'd3326,  18'd1794,  18'd3853,  -18'd2464,  -18'd2613,  18'd3573,  -18'd7681,  -18'd4782,  18'd4181,  18'd7636,  18'd1946,  -18'd9321,  -18'd33,  
-18'd1596,  -18'd3491,  18'd5463,  -18'd4080,  18'd8567,  -18'd8537,  18'd3232,  -18'd8366,  -18'd8699,  18'd5873,  -18'd9441,  -18'd12127,  18'd6608,  -18'd8845,  18'd1920,  18'd8420,  
-18'd4936,  -18'd647,  -18'd3544,  -18'd426,  -18'd8482,  18'd7195,  -18'd644,  18'd1126,  -18'd9979,  -18'd14343,  18'd2262,  -18'd2744,  18'd511,  -18'd4165,  18'd2593,  -18'd9673,  

18'd4967,  18'd20907,  18'd5608,  18'd14038,  18'd8798,  18'd2783,  18'd9264,  -18'd1639,  -18'd5929,  -18'd14643,  -18'd1165,  -18'd22979,  18'd9588,  -18'd7526,  18'd1238,  18'd17943,  
-18'd4472,  -18'd10470,  18'd8183,  -18'd312,  18'd5297,  -18'd14112,  18'd10408,  18'd4653,  -18'd21973,  -18'd1473,  18'd16349,  -18'd8339,  18'd276,  -18'd5371,  18'd13328,  -18'd9759,  
-18'd15599,  18'd9817,  18'd12034,  -18'd9,  -18'd8943,  -18'd1766,  -18'd4058,  18'd16982,  18'd2721,  18'd2286,  18'd9211,  18'd3066,  -18'd5495,  18'd7699,  -18'd4821,  18'd725,  
-18'd10756,  18'd24011,  -18'd1577,  -18'd2903,  -18'd3488,  -18'd6882,  18'd5648,  18'd12434,  -18'd7215,  -18'd8516,  -18'd14152,  18'd14224,  -18'd1318,  -18'd470,  18'd2145,  -18'd15304,  
-18'd5449,  -18'd5745,  18'd762,  18'd31876,  18'd8191,  18'd8541,  18'd4341,  -18'd1888,  18'd7895,  18'd3170,  -18'd1174,  18'd1120,  18'd6436,  18'd4383,  -18'd3734,  18'd13321,  
-18'd6690,  18'd6437,  -18'd2188,  -18'd5408,  18'd1583,  -18'd4587,  -18'd13807,  18'd13583,  -18'd22186,  18'd8383,  18'd9644,  18'd5424,  18'd666,  18'd796,  18'd1631,  18'd3616,  
-18'd7894,  18'd24166,  18'd968,  -18'd9570,  -18'd3937,  18'd11170,  -18'd25139,  18'd1495,  -18'd7599,  -18'd4179,  18'd4109,  18'd1138,  18'd7759,  18'd17111,  18'd2486,  18'd19475,  
-18'd16866,  18'd28120,  18'd2984,  -18'd5038,  -18'd7304,  -18'd5292,  -18'd26196,  18'd2469,  -18'd7506,  18'd5590,  -18'd12863,  18'd4057,  18'd2346,  18'd2512,  -18'd1789,  18'd16031,  
18'd10487,  -18'd1652,  18'd1764,  -18'd25236,  -18'd9441,  18'd5273,  18'd3355,  -18'd2614,  18'd7111,  -18'd15036,  -18'd8215,  -18'd10680,  18'd3119,  18'd10285,  -18'd4737,  18'd2192,  
18'd11556,  -18'd10677,  -18'd5149,  18'd13998,  18'd536,  -18'd11392,  -18'd23779,  18'd10396,  18'd4611,  -18'd2405,  -18'd9035,  -18'd898,  18'd2621,  18'd5351,  -18'd1300,  -18'd966,  
18'd2422,  18'd7102,  -18'd3176,  -18'd4613,  18'd2305,  -18'd6249,  -18'd3882,  18'd11325,  18'd456,  18'd13786,  18'd8349,  18'd6461,  18'd2837,  18'd150,  18'd4257,  -18'd2122,  
18'd2471,  18'd5899,  -18'd15,  18'd6059,  18'd0,  -18'd5255,  -18'd21766,  -18'd12437,  -18'd3185,  18'd19774,  18'd8773,  18'd11989,  -18'd4947,  18'd6860,  18'd6546,  18'd27496,  
-18'd3851,  18'd17951,  18'd8297,  -18'd13286,  -18'd3944,  18'd2778,  18'd7394,  18'd9680,  18'd1334,  -18'd1892,  18'd7060,  -18'd12756,  -18'd8055,  18'd5833,  -18'd493,  18'd7713,  
-18'd1249,  18'd9100,  18'd8785,  18'd16838,  18'd5296,  -18'd19245,  -18'd24217,  18'd81,  -18'd3959,  -18'd17789,  18'd3736,  -18'd13752,  18'd2325,  18'd169,  -18'd5306,  18'd6302,  
-18'd12736,  18'd10507,  18'd542,  18'd674,  -18'd2034,  -18'd11901,  -18'd13520,  -18'd2778,  -18'd12295,  18'd2415,  -18'd3413,  -18'd6549,  -18'd2567,  -18'd7915,  18'd7758,  -18'd9421,  
-18'd7271,  -18'd5461,  -18'd15650,  18'd7471,  -18'd5164,  -18'd5173,  -18'd1561,  -18'd743,  -18'd5276,  -18'd1990,  -18'd2087,  18'd273,  18'd9518,  -18'd4313,  18'd14725,  -18'd8973,  

-18'd341,  -18'd4005,  -18'd3295,  18'd1066,  18'd8686,  18'd3124,  -18'd829,  -18'd6525,  -18'd7255,  18'd5212,  18'd1778,  -18'd5740,  -18'd7689,  -18'd7556,  18'd3558,  -18'd12625,  
-18'd7936,  -18'd762,  -18'd859,  18'd3127,  18'd8867,  -18'd11109,  -18'd8856,  -18'd4574,  -18'd9549,  18'd3215,  -18'd5117,  -18'd11209,  -18'd4444,  -18'd179,  -18'd1336,  -18'd9705,  
-18'd10458,  -18'd5197,  18'd2726,  18'd569,  18'd5545,  -18'd2102,  -18'd4395,  -18'd7738,  -18'd6546,  18'd370,  -18'd6966,  -18'd5154,  18'd1870,  -18'd6012,  -18'd2259,  -18'd13320,  
-18'd5080,  18'd14,  -18'd8989,  -18'd10706,  18'd5805,  -18'd6218,  -18'd12924,  -18'd3104,  -18'd7994,  18'd4907,  18'd23,  -18'd5179,  18'd2264,  18'd3026,  18'd1883,  -18'd1885,  
-18'd4341,  -18'd2968,  -18'd213,  -18'd7352,  18'd7107,  -18'd1454,  -18'd9434,  -18'd4881,  18'd4009,  -18'd9690,  -18'd6557,  -18'd2655,  -18'd2666,  18'd1563,  18'd2720,  18'd685,  
-18'd5665,  -18'd6214,  -18'd13961,  18'd844,  18'd6402,  -18'd2932,  -18'd1440,  -18'd8636,  18'd1302,  18'd3957,  -18'd1433,  -18'd13465,  18'd1333,  -18'd11559,  -18'd7958,  -18'd755,  
18'd2591,  -18'd11375,  18'd1740,  -18'd14107,  -18'd4802,  -18'd8551,  -18'd1402,  -18'd5328,  -18'd9629,  18'd377,  18'd4852,  18'd2963,  18'd2555,  -18'd9649,  -18'd12087,  -18'd11977,  
-18'd9817,  18'd342,  -18'd10801,  18'd4699,  18'd8880,  -18'd11724,  -18'd3913,  -18'd8075,  18'd2097,  -18'd8351,  -18'd9349,  -18'd11700,  18'd4938,  -18'd11433,  18'd1385,  18'd778,  
18'd1570,  -18'd10025,  -18'd5031,  18'd6567,  18'd5797,  18'd2426,  -18'd9060,  18'd3592,  -18'd1338,  18'd3920,  -18'd8165,  -18'd6869,  18'd5544,  -18'd5798,  18'd2973,  18'd3123,  
-18'd4624,  18'd1551,  -18'd7493,  -18'd5368,  -18'd3196,  -18'd11270,  18'd246,  -18'd5318,  -18'd5165,  18'd1256,  18'd664,  18'd1778,  18'd471,  18'd5378,  -18'd4107,  -18'd11323,  
-18'd7584,  18'd3381,  -18'd6553,  18'd1875,  18'd8682,  -18'd1733,  18'd1593,  18'd6534,  18'd2676,  18'd4918,  -18'd7522,  18'd2419,  -18'd2829,  18'd5700,  -18'd8845,  -18'd6322,  
-18'd317,  -18'd4790,  -18'd7521,  18'd2185,  -18'd7640,  -18'd3088,  -18'd335,  -18'd7460,  -18'd9364,  -18'd10243,  -18'd10643,  -18'd1624,  18'd4282,  18'd3867,  -18'd8690,  -18'd1466,  
-18'd10189,  -18'd7574,  -18'd7302,  18'd3192,  18'd8448,  18'd3548,  -18'd6027,  18'd3993,  -18'd4266,  18'd4941,  -18'd9330,  -18'd11278,  18'd7648,  18'd2613,  -18'd4312,  -18'd6552,  
-18'd11611,  18'd3892,  18'd4320,  18'd6597,  -18'd627,  -18'd15,  -18'd8773,  -18'd2893,  -18'd2225,  18'd6923,  -18'd2038,  18'd2769,  -18'd6062,  18'd4725,  18'd402,  -18'd1448,  
-18'd3687,  -18'd11241,  -18'd9799,  -18'd6281,  18'd6065,  18'd1295,  -18'd9826,  -18'd3781,  -18'd2316,  18'd4629,  18'd5097,  -18'd5325,  -18'd2374,  -18'd99,  18'd5869,  -18'd30,  
-18'd1524,  -18'd7454,  -18'd1653,  -18'd5194,  -18'd3941,  -18'd6987,  -18'd4320,  18'd4034,  18'd1177,  18'd3317,  18'd2763,  18'd1376,  -18'd7183,  -18'd11799,  -18'd733,  18'd545,  

18'd8291,  -18'd17975,  -18'd16398,  18'd819,  18'd1560,  18'd4790,  -18'd2097,  18'd828,  18'd19477,  -18'd9283,  -18'd13841,  18'd3190,  -18'd5661,  18'd3045,  -18'd4745,  -18'd13383,  
18'd24414,  -18'd3481,  -18'd9638,  18'd2073,  18'd7975,  18'd7494,  18'd17968,  -18'd12065,  18'd7527,  18'd15909,  18'd2207,  18'd10500,  -18'd963,  18'd1107,  18'd2826,  -18'd16089,  
18'd15960,  -18'd2910,  18'd15195,  -18'd3489,  -18'd4023,  -18'd15482,  18'd14787,  -18'd2216,  18'd12771,  18'd15599,  -18'd3277,  18'd21409,  18'd6315,  -18'd601,  18'd8670,  -18'd4817,  
-18'd3488,  18'd17827,  18'd23976,  -18'd19184,  18'd924,  -18'd14133,  18'd19926,  18'd13805,  18'd464,  -18'd488,  18'd854,  18'd13564,  18'd4116,  18'd2669,  -18'd1337,  -18'd1380,  
-18'd6803,  18'd6730,  -18'd2201,  18'd15588,  18'd8305,  18'd11399,  18'd1695,  18'd637,  18'd12075,  18'd1152,  18'd2290,  18'd1412,  18'd8197,  18'd4001,  -18'd10,  18'd16215,  
18'd7368,  -18'd9765,  -18'd10706,  18'd17873,  18'd4845,  18'd3633,  18'd9131,  -18'd3627,  -18'd1816,  18'd16163,  -18'd3081,  18'd5380,  -18'd3401,  18'd6398,  -18'd11004,  18'd679,  
-18'd9570,  18'd3385,  -18'd11952,  18'd5681,  -18'd5991,  -18'd6195,  -18'd6609,  18'd700,  18'd5193,  18'd25131,  18'd4372,  18'd26703,  18'd8742,  -18'd2388,  -18'd4,  -18'd9438,  
-18'd12751,  18'd2743,  18'd1604,  -18'd7980,  18'd2231,  18'd1743,  -18'd3753,  18'd5549,  -18'd11257,  -18'd3262,  18'd33549,  18'd19331,  -18'd4546,  18'd9343,  18'd10429,  18'd582,  
-18'd12027,  -18'd17218,  -18'd94,  -18'd18767,  -18'd7952,  -18'd1393,  18'd13342,  -18'd3318,  -18'd735,  18'd3053,  -18'd1191,  -18'd3219,  -18'd939,  -18'd6875,  18'd7892,  18'd4182,  
18'd7705,  -18'd8413,  -18'd1314,  18'd1,  -18'd2816,  18'd1339,  18'd9797,  -18'd11194,  18'd2059,  18'd5091,  18'd16911,  -18'd699,  -18'd1843,  -18'd4048,  -18'd1268,  18'd13126,  
-18'd8308,  -18'd4893,  -18'd17743,  18'd5060,  18'd8713,  -18'd7622,  -18'd19309,  18'd7885,  -18'd5813,  18'd19291,  18'd4576,  18'd16197,  18'd7718,  -18'd4697,  18'd2629,  -18'd3238,  
-18'd11474,  -18'd28395,  -18'd5075,  -18'd5083,  18'd5761,  -18'd22390,  -18'd2188,  18'd13628,  -18'd8648,  -18'd3923,  18'd19969,  18'd13691,  -18'd5739,  18'd2042,  -18'd4051,  -18'd12217,  
-18'd1376,  -18'd419,  18'd10452,  -18'd21365,  -18'd5003,  18'd6639,  18'd17855,  18'd11511,  18'd8163,  -18'd3261,  18'd12371,  -18'd6083,  -18'd4675,  -18'd9880,  18'd13816,  -18'd13610,  
18'd3733,  -18'd14366,  18'd16270,  -18'd15144,  18'd6182,  18'd1561,  18'd11021,  18'd22114,  18'd4411,  18'd10316,  18'd1643,  -18'd1577,  18'd7931,  -18'd12648,  -18'd12515,  18'd1342,  
18'd10635,  -18'd7382,  -18'd9586,  18'd717,  -18'd7774,  18'd1000,  18'd1783,  -18'd12450,  -18'd4561,  -18'd2082,  18'd4034,  18'd6494,  -18'd6688,  18'd4057,  -18'd250,  18'd5257,  
18'd15519,  -18'd6123,  -18'd15433,  18'd3696,  -18'd4312,  -18'd16078,  -18'd8382,  18'd9479,  18'd2644,  18'd14479,  18'd3493,  18'd8378,  18'd3756,  18'd2335,  18'd4722,  -18'd12991,  

18'd26887,  -18'd6883,  18'd11150,  18'd7037,  18'd5948,  18'd6634,  18'd13272,  -18'd4547,  18'd18845,  18'd16876,  18'd9479,  18'd14992,  18'd1067,  18'd5803,  18'd14862,  18'd8739,  
18'd4730,  -18'd2630,  -18'd6334,  18'd27842,  18'd3758,  18'd5617,  18'd7222,  -18'd903,  18'd20038,  18'd3437,  18'd8109,  18'd17843,  -18'd10462,  18'd11735,  18'd3079,  18'd12900,  
-18'd12678,  18'd16304,  18'd10570,  18'd6684,  -18'd7535,  -18'd6655,  -18'd9680,  18'd5542,  18'd1649,  -18'd20076,  18'd930,  -18'd1652,  18'd7762,  18'd9401,  -18'd28726,  18'd7694,  
-18'd18568,  18'd22467,  18'd6384,  18'd11122,  -18'd3286,  18'd19493,  -18'd18784,  18'd4459,  -18'd12736,  -18'd3405,  -18'd14499,  18'd10315,  -18'd7836,  18'd10136,  -18'd4253,  -18'd690,  
18'd13564,  -18'd8820,  -18'd7464,  -18'd6533,  -18'd144,  18'd429,  18'd3698,  18'd3291,  -18'd3614,  -18'd13055,  -18'd4640,  18'd9682,  18'd5473,  18'd8263,  18'd4925,  -18'd8767,  
-18'd5799,  18'd2693,  -18'd5047,  -18'd14471,  -18'd5262,  -18'd1538,  -18'd5816,  -18'd1971,  -18'd3749,  -18'd5285,  18'd22485,  18'd27619,  -18'd1346,  18'd7865,  18'd19818,  18'd449,  
18'd5431,  -18'd4410,  18'd13333,  -18'd13770,  -18'd1808,  18'd1234,  -18'd13664,  -18'd14366,  18'd10274,  18'd56,  18'd220,  18'd344,  -18'd5628,  18'd9835,  -18'd11912,  18'd6545,  
18'd10464,  18'd29836,  -18'd11697,  18'd12843,  -18'd1923,  18'd68,  -18'd28128,  -18'd15094,  -18'd1244,  18'd18159,  -18'd17390,  18'd11860,  18'd7484,  18'd10428,  -18'd4681,  18'd10033,  
18'd4337,  18'd8109,  18'd10151,  -18'd11001,  18'd6607,  -18'd1715,  -18'd13171,  -18'd1528,  -18'd3678,  -18'd17522,  -18'd656,  -18'd8151,  18'd7469,  -18'd374,  18'd1384,  18'd5531,  
-18'd4400,  18'd569,  18'd1193,  -18'd21707,  18'd3108,  -18'd16827,  -18'd8855,  18'd12440,  18'd543,  -18'd5762,  18'd3158,  18'd382,  -18'd3733,  -18'd3494,  -18'd775,  -18'd161,  
18'd10407,  18'd9007,  18'd11993,  -18'd5164,  -18'd8993,  -18'd3334,  18'd18603,  -18'd3953,  18'd5092,  -18'd1277,  18'd898,  -18'd9093,  18'd5946,  -18'd11941,  18'd1693,  -18'd3847,  
18'd7461,  18'd30283,  -18'd13695,  -18'd1892,  18'd8657,  18'd8856,  18'd9764,  18'd7487,  18'd4834,  18'd8393,  -18'd8678,  18'd4900,  18'd7840,  18'd1918,  18'd4387,  18'd19842,  
18'd4957,  18'd15383,  -18'd2345,  -18'd6337,  18'd5181,  -18'd6735,  -18'd2611,  18'd6629,  -18'd2643,  -18'd6900,  18'd6644,  -18'd18291,  -18'd8046,  -18'd13797,  18'd3624,  18'd26067,  
18'd5683,  18'd4434,  -18'd3500,  -18'd518,  -18'd2251,  -18'd17816,  -18'd722,  18'd5134,  -18'd2900,  18'd17380,  18'd1991,  -18'd11458,  -18'd7634,  -18'd8092,  18'd9713,  18'd7384,  
-18'd657,  -18'd16760,  18'd7629,  -18'd6149,  -18'd1963,  18'd218,  18'd9731,  18'd1627,  -18'd806,  18'd8062,  -18'd10132,  -18'd8520,  18'd3398,  -18'd9924,  18'd5011,  -18'd6088,  
-18'd20060,  18'd1482,  -18'd3842,  18'd14808,  18'd6967,  -18'd10289,  18'd11419,  18'd13947,  18'd1409,  -18'd1867,  18'd1452,  -18'd13248,  -18'd7852,  -18'd14947,  18'd5031,  18'd8583,  

18'd12510,  -18'd26631,  -18'd9082,  18'd626,  18'd6550,  18'd4357,  -18'd1774,  -18'd8648,  18'd13907,  18'd21680,  -18'd21100,  18'd31247,  18'd3192,  18'd38521,  -18'd5851,  18'd7365,  
18'd5985,  -18'd23314,  -18'd20043,  18'd24288,  -18'd4232,  -18'd27425,  -18'd11571,  -18'd14969,  -18'd9160,  18'd18002,  -18'd7542,  18'd3370,  18'd6128,  18'd3561,  18'd6725,  -18'd8364,  
18'd10643,  -18'd27539,  -18'd2862,  18'd11202,  -18'd1014,  -18'd7097,  18'd23411,  -18'd5858,  -18'd30356,  18'd16845,  18'd12036,  -18'd605,  -18'd6103,  18'd1256,  18'd12657,  -18'd16796,  
18'd11325,  -18'd21451,  18'd9872,  -18'd2366,  -18'd3596,  18'd10296,  18'd293,  18'd2582,  18'd11895,  -18'd2706,  18'd6141,  18'd4635,  -18'd3529,  18'd9781,  18'd10014,  -18'd5941,  
18'd17314,  18'd3709,  18'd4912,  18'd23605,  -18'd4845,  -18'd487,  -18'd1466,  -18'd6812,  -18'd4877,  18'd1268,  -18'd9718,  18'd1371,  18'd10415,  -18'd1789,  18'd3651,  -18'd11614,  
18'd6093,  -18'd2839,  -18'd14160,  18'd21590,  -18'd683,  -18'd8491,  18'd448,  18'd2559,  -18'd4198,  18'd3909,  -18'd2594,  -18'd10192,  18'd9565,  18'd2397,  18'd9400,  -18'd1169,  
18'd2140,  18'd879,  -18'd5873,  -18'd7416,  -18'd555,  18'd5516,  18'd24525,  -18'd5454,  -18'd2543,  18'd3814,  18'd11316,  18'd9105,  18'd2891,  -18'd890,  18'd1430,  -18'd8513,  
18'd6523,  18'd7386,  18'd8865,  -18'd15653,  -18'd3274,  18'd1459,  18'd4667,  -18'd4152,  18'd25145,  18'd13438,  18'd1962,  18'd13043,  18'd9584,  18'd10963,  18'd752,  18'd6108,  
-18'd9460,  18'd10323,  18'd7772,  18'd4509,  18'd6448,  18'd763,  -18'd1632,  18'd10218,  -18'd2644,  18'd13107,  18'd547,  18'd1142,  -18'd532,  -18'd3129,  18'd1329,  18'd13125,  
-18'd187,  18'd2283,  -18'd925,  18'd5446,  -18'd1983,  -18'd4080,  18'd7200,  -18'd4824,  -18'd9897,  18'd1314,  -18'd3628,  -18'd15038,  -18'd2488,  -18'd433,  18'd14395,  -18'd51,  
-18'd4974,  -18'd9828,  18'd1356,  -18'd16531,  -18'd7304,  18'd21673,  18'd11884,  18'd8790,  18'd4235,  -18'd10478,  18'd6792,  18'd2305,  -18'd4098,  18'd1169,  -18'd2288,  -18'd13142,  
-18'd1495,  -18'd5961,  18'd4330,  -18'd4236,  -18'd6244,  18'd3336,  -18'd5735,  18'd1870,  18'd16654,  18'd6325,  -18'd1316,  18'd7429,  18'd4111,  -18'd2695,  18'd1763,  18'd6176,  
-18'd9674,  -18'd7467,  18'd12870,  18'd17358,  -18'd5515,  18'd1957,  18'd7715,  -18'd5339,  18'd4231,  18'd5256,  18'd1087,  18'd10533,  -18'd2683,  -18'd4590,  18'd12497,  18'd14181,  
18'd40,  -18'd8328,  -18'd3854,  -18'd236,  -18'd5360,  18'd8217,  18'd12247,  -18'd8838,  -18'd11341,  -18'd7459,  18'd5476,  18'd7577,  18'd5257,  18'd3853,  18'd14791,  -18'd656,  
-18'd5193,  18'd5919,  18'd6736,  -18'd340,  -18'd5784,  18'd7168,  18'd23675,  18'd8903,  18'd4575,  18'd8073,  18'd10407,  -18'd5957,  18'd1176,  18'd1332,  18'd6945,  18'd3826,  
-18'd5752,  -18'd9400,  -18'd17531,  18'd8169,  -18'd8188,  18'd2702,  -18'd586,  -18'd7691,  -18'd3949,  18'd1784,  -18'd7665,  -18'd7618,  18'd4096,  18'd9036,  18'd6977,  18'd9908,  

18'd13226,  -18'd4652,  -18'd2106,  18'd32237,  18'd6906,  -18'd8880,  18'd2846,  -18'd4273,  -18'd2643,  18'd628,  18'd15962,  -18'd3298,  -18'd2087,  -18'd2261,  -18'd4283,  18'd31872,  
-18'd7516,  -18'd13471,  -18'd2999,  -18'd5861,  18'd368,  18'd6472,  18'd13378,  -18'd4437,  18'd17249,  18'd16927,  18'd9549,  18'd16232,  -18'd7813,  18'd3873,  -18'd5642,  18'd1914,  
18'd10630,  -18'd14065,  -18'd7318,  18'd20892,  18'd2192,  18'd5745,  -18'd9839,  -18'd12915,  18'd13664,  -18'd19750,  -18'd25482,  -18'd16544,  18'd6612,  18'd6964,  -18'd23592,  -18'd1054,  
18'd32,  -18'd23204,  -18'd16474,  -18'd9568,  -18'd2498,  18'd8477,  18'd16374,  -18'd2793,  -18'd21821,  18'd11490,  18'd3976,  -18'd11317,  -18'd7907,  -18'd1522,  -18'd2911,  -18'd9219,  
-18'd5633,  -18'd12634,  18'd4873,  18'd27384,  -18'd7778,  -18'd13797,  18'd2650,  18'd2065,  -18'd5447,  18'd5308,  -18'd8748,  18'd1480,  -18'd5643,  18'd3736,  -18'd9999,  -18'd5549,  
18'd2117,  -18'd2465,  18'd2990,  -18'd6690,  18'd6716,  18'd5978,  -18'd303,  18'd1509,  -18'd8652,  -18'd1433,  18'd2094,  18'd645,  -18'd5909,  18'd11281,  -18'd682,  18'd1976,  
-18'd3650,  -18'd17523,  -18'd14094,  18'd10646,  -18'd4318,  -18'd7257,  -18'd12474,  -18'd15964,  18'd14701,  18'd16259,  18'd13469,  18'd5164,  18'd2795,  18'd9571,  18'd5771,  -18'd21348,  
18'd7933,  18'd305,  -18'd18805,  -18'd4468,  -18'd4159,  18'd9712,  -18'd3492,  18'd8472,  -18'd8561,  -18'd15804,  18'd10265,  18'd1336,  -18'd7564,  -18'd1717,  18'd10484,  -18'd19071,  
18'd2674,  -18'd23015,  18'd404,  18'd9494,  -18'd4690,  -18'd2635,  18'd5681,  -18'd12043,  -18'd3182,  18'd19107,  -18'd12118,  18'd1660,  18'd5441,  18'd7729,  -18'd10252,  -18'd6502,  
18'd6654,  -18'd9827,  18'd4753,  -18'd6824,  -18'd7207,  -18'd26102,  -18'd8938,  -18'd3157,  -18'd5842,  -18'd7850,  18'd5263,  18'd4930,  18'd5594,  -18'd1227,  18'd2050,  -18'd4996,  
18'd7987,  -18'd7202,  18'd4087,  -18'd4193,  18'd6951,  18'd12719,  18'd6634,  -18'd613,  18'd3417,  18'd14252,  -18'd137,  -18'd6770,  -18'd712,  18'd12442,  18'd373,  -18'd12163,  
18'd8256,  -18'd16773,  -18'd17355,  18'd1603,  -18'd5040,  -18'd10083,  18'd6785,  -18'd5644,  18'd6541,  -18'd20876,  -18'd824,  -18'd8670,  -18'd3771,  -18'd20111,  18'd19735,  18'd8859,  
-18'd285,  -18'd9656,  18'd2288,  18'd6344,  18'd5761,  18'd9548,  18'd2883,  -18'd9818,  -18'd3625,  18'd72,  18'd11765,  18'd6556,  18'd7357,  18'd12185,  -18'd11841,  18'd9414,  
18'd8092,  -18'd13997,  18'd2069,  -18'd10493,  -18'd7303,  18'd3892,  18'd8347,  -18'd587,  -18'd3850,  18'd12509,  18'd10723,  18'd17096,  -18'd5684,  -18'd116,  18'd5986,  18'd11377,  
18'd19482,  18'd4683,  18'd1237,  18'd3524,  18'd3161,  18'd21520,  18'd35608,  -18'd324,  18'd11926,  18'd4424,  -18'd95,  18'd2845,  -18'd3873,  -18'd7451,  18'd6466,  18'd3901,  
18'd2545,  -18'd4674,  18'd3283,  18'd3847,  -18'd495,  -18'd6129,  18'd18892,  -18'd15533,  18'd12703,  -18'd19368,  -18'd3724,  -18'd19881,  18'd6176,  -18'd14732,  18'd6856,  18'd3818,  

18'd14055,  18'd23622,  18'd2730,  -18'd17865,  -18'd8202,  18'd3555,  -18'd10879,  18'd6371,  18'd7493,  18'd11048,  -18'd1545,  18'd19554,  -18'd3687,  -18'd683,  -18'd4823,  -18'd9539,  
18'd7618,  18'd11354,  18'd2081,  18'd7210,  18'd5114,  18'd9393,  -18'd905,  -18'd4860,  18'd19781,  -18'd5808,  18'd4826,  18'd9612,  -18'd5295,  -18'd527,  -18'd10835,  -18'd3250,  
18'd16027,  18'd3352,  -18'd9167,  18'd300,  18'd2643,  -18'd5777,  18'd7793,  -18'd4593,  18'd7401,  18'd3181,  -18'd16542,  18'd4226,  -18'd3282,  -18'd7796,  -18'd5407,  -18'd1483,  
-18'd4440,  -18'd3981,  18'd7060,  18'd12161,  18'd7399,  -18'd1493,  18'd27519,  -18'd1156,  -18'd3906,  18'd122,  18'd770,  18'd305,  -18'd5545,  18'd3981,  -18'd7151,  -18'd12346,  
18'd12353,  18'd27771,  18'd9674,  -18'd15129,  18'd4707,  -18'd8837,  -18'd5628,  18'd13814,  18'd4026,  18'd14695,  -18'd7420,  18'd11330,  -18'd9601,  18'd12999,  18'd3098,  18'd17262,  
-18'd20412,  18'd4174,  18'd595,  18'd17196,  18'd7803,  18'd9507,  -18'd1074,  -18'd8850,  18'd17279,  18'd19912,  -18'd7639,  18'd4221,  -18'd2284,  18'd7950,  -18'd9157,  18'd14871,  
18'd6430,  -18'd15974,  -18'd1292,  18'd5413,  18'd5563,  18'd8359,  18'd4301,  18'd6947,  18'd7059,  -18'd14341,  18'd4121,  -18'd1740,  -18'd6832,  -18'd13178,  -18'd4145,  18'd4276,  
-18'd2301,  -18'd22814,  18'd20312,  -18'd10627,  18'd5325,  18'd20395,  18'd29182,  -18'd10943,  18'd9379,  -18'd15678,  18'd18399,  -18'd5420,  18'd2475,  -18'd577,  18'd16939,  -18'd33561,  
18'd9483,  18'd5430,  -18'd318,  18'd15508,  18'd7629,  -18'd9993,  -18'd16575,  18'd5029,  18'd4087,  18'd15963,  18'd5544,  18'd7489,  -18'd743,  18'd4020,  18'd4031,  18'd4994,  
18'd5215,  -18'd624,  -18'd1823,  -18'd5052,  -18'd404,  -18'd8293,  -18'd19374,  -18'd5518,  -18'd2611,  18'd13576,  -18'd1173,  18'd7097,  18'd1039,  18'd10462,  18'd13190,  -18'd781,  
18'd5232,  -18'd1185,  18'd3373,  18'd3763,  18'd6353,  -18'd9190,  -18'd16567,  18'd16270,  -18'd13682,  -18'd7483,  18'd8510,  -18'd7615,  18'd6608,  -18'd10149,  18'd7452,  18'd1656,  
-18'd5154,  18'd30797,  18'd3532,  -18'd1986,  -18'd7983,  18'd14771,  18'd17541,  18'd34327,  18'd7014,  -18'd12047,  18'd2666,  -18'd9366,  -18'd3196,  -18'd15213,  -18'd12084,  -18'd774,  
18'd26624,  18'd7451,  -18'd10615,  -18'd5505,  18'd2822,  -18'd6577,  -18'd15972,  -18'd12181,  18'd9240,  18'd15091,  -18'd1132,  18'd52,  18'd7045,  18'd3885,  -18'd13163,  18'd10542,  
18'd12642,  -18'd10610,  -18'd373,  18'd3875,  -18'd7974,  -18'd16706,  -18'd920,  18'd15482,  18'd6943,  18'd3293,  -18'd2500,  -18'd142,  -18'd1744,  18'd1553,  18'd7171,  -18'd5815,  
-18'd6422,  -18'd7860,  -18'd7196,  18'd1126,  18'd4984,  -18'd28313,  -18'd5307,  18'd13737,  -18'd7916,  -18'd587,  18'd524,  -18'd14983,  18'd1305,  18'd2545,  18'd4229,  -18'd4954,  
-18'd995,  18'd2364,  18'd5806,  -18'd1527,  -18'd8014,  -18'd5695,  18'd8769,  18'd21204,  18'd2400,  18'd6471,  -18'd5307,  18'd1747,  18'd2171,  -18'd2046,  18'd2938,  -18'd4005,  

-18'd155,  18'd6459,  18'd10836,  18'd17373,  -18'd7454,  -18'd13973,  -18'd2686,  18'd9312,  -18'd6074,  18'd4332,  18'd2030,  -18'd20466,  18'd7759,  18'd4398,  -18'd122,  18'd9861,  
18'd4907,  18'd18654,  18'd12095,  -18'd16633,  18'd7943,  18'd12614,  18'd8361,  18'd55,  18'd6917,  18'd4891,  18'd12403,  -18'd4528,  -18'd3816,  18'd6587,  18'd799,  18'd13113,  
18'd2199,  18'd12728,  18'd833,  -18'd6650,  -18'd47,  18'd8053,  -18'd3190,  18'd6017,  18'd20134,  18'd2855,  -18'd8774,  18'd14182,  18'd1852,  18'd19345,  -18'd1245,  18'd16079,  
-18'd9445,  18'd4920,  -18'd2798,  18'd8629,  -18'd1188,  -18'd13341,  18'd9337,  -18'd16701,  -18'd5881,  18'd8959,  18'd311,  -18'd1277,  18'd1050,  -18'd5790,  -18'd336,  18'd4501,  
-18'd14459,  -18'd1986,  18'd3644,  18'd22419,  18'd5859,  18'd14062,  -18'd8351,  18'd2714,  18'd3407,  18'd23994,  -18'd5705,  18'd21177,  18'd1363,  18'd8113,  18'd2632,  -18'd1885,  
-18'd5037,  18'd7685,  18'd6077,  -18'd3775,  18'd6411,  18'd19798,  -18'd8235,  -18'd6166,  18'd7189,  -18'd6800,  -18'd757,  18'd9034,  18'd4438,  18'd16123,  -18'd17810,  18'd12959,  
18'd1777,  18'd6757,  -18'd6585,  18'd11159,  18'd1493,  -18'd5326,  -18'd33653,  -18'd754,  18'd6285,  18'd5675,  -18'd12141,  18'd2741,  -18'd2750,  18'd16450,  18'd7225,  18'd9117,  
-18'd9973,  -18'd2949,  -18'd22259,  18'd8552,  18'd940,  -18'd20247,  -18'd17676,  18'd4098,  18'd1673,  18'd12227,  -18'd5689,  18'd11387,  -18'd1295,  18'd6233,  -18'd2871,  18'd126,  
18'd9617,  -18'd17824,  -18'd5525,  -18'd19841,  -18'd249,  -18'd319,  -18'd6396,  -18'd15771,  18'd5892,  18'd8336,  18'd1705,  18'd1041,  -18'd1499,  -18'd2864,  18'd204,  -18'd11670,  
18'd13284,  -18'd2638,  -18'd5085,  -18'd8787,  18'd7009,  18'd4667,  -18'd6354,  18'd5685,  18'd5688,  -18'd16531,  18'd3896,  -18'd9444,  18'd9544,  18'd685,  18'd564,  -18'd5156,  
18'd4341,  -18'd8349,  -18'd10568,  -18'd11607,  18'd2383,  -18'd7749,  -18'd2016,  -18'd17565,  -18'd12952,  18'd6795,  18'd1361,  -18'd5259,  -18'd5796,  -18'd7430,  18'd11290,  18'd11005,  
-18'd4193,  -18'd2356,  -18'd20314,  18'd11383,  -18'd7834,  -18'd12818,  -18'd8502,  -18'd5212,  18'd4519,  18'd4044,  18'd529,  18'd6312,  18'd3146,  -18'd3002,  18'd8370,  -18'd1840,  
18'd15603,  18'd7920,  18'd7669,  -18'd29612,  -18'd4507,  -18'd3193,  18'd1503,  18'd9355,  18'd3497,  -18'd3551,  18'd2223,  18'd11,  18'd1198,  -18'd5738,  18'd2795,  -18'd15962,  
-18'd10331,  18'd758,  18'd1104,  18'd3287,  -18'd5703,  -18'd12046,  18'd11234,  18'd1491,  18'd5360,  -18'd23628,  18'd12647,  -18'd12703,  -18'd3155,  -18'd5523,  -18'd3565,  18'd883,  
-18'd570,  -18'd1242,  -18'd5836,  18'd3537,  18'd5027,  -18'd5886,  18'd1758,  -18'd7121,  -18'd16782,  18'd2677,  -18'd8868,  -18'd15613,  18'd1036,  -18'd14625,  18'd4121,  -18'd10662,  
-18'd2550,  -18'd10376,  18'd1949,  -18'd2853,  18'd1085,  18'd3717,  18'd2737,  -18'd5965,  18'd3933,  18'd13173,  18'd7214,  -18'd5672,  18'd5814,  -18'd12109,  18'd7637,  -18'd23355
	};
	
	always @(posedge clk) begin
		if (rstn == 0) begin
			qa <= 0;
		end
		else if (!cena) begin
			qa <= weight[aa];
		end
	end
	
endmodule




