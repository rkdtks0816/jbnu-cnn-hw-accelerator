 `include "global.sv"
`include "timescale.sv"

module sign_mnist(
	input			clk,
	input			rstn,
	input			en,
	input				key_1,
	
	output	reg				ready,
	output			[`WD:0]	q_data,
	output	reg				push
	);
	reg	[`WD:0]		dt;
	
	reg	[1:0]		din;
	
	reg	[4:0]		count;
	
	reg	[10:0]		cnt;
	reg					cnt_en;
	wire			cnt_max = cnt == 10'd783;
	wire			end_cnt_en = cnt_max;
	

	always @(posedge clk, negedge rstn) begin
		if(rstn == 0) begin
			din	<=	2'd0;
			push	<=	1'b0;
		end
		else begin
			if(en == 1) begin
				din[0]	<=	key_1;
				din[1]	<=	din[0];
				if(din[0] == 1 && din[1] == 0) begin
					push	<=	1'b1;
				end
				else begin
					push	<=	1'b0;
				end
			end
			else begin
				din	<=	2'b0;
				push	<=	1'b0;
			end
		end
	end

	always @(posedge clk, negedge rstn) begin
		if (rstn == 0) begin
			count	<=	5'd31;
		end
		else begin
			if(en == 1) begin
				if(push == 1) begin
					count	<=	count + 1;
				end
			end
			else begin
				count	<=	5'd31;
			end
		end
	end

	always @(posedge clk)
		if (`RST)			cnt_en <= 0;
		else if (push)			cnt_en <= 1;
		else if (end_cnt_en)		cnt_en <= 0;

	always @(posedge clk)
		if (`RST)	cnt <= 0;
		else if(cnt_en)	cnt <= cnt_max? 0: cnt + 1;

	always @(posedge clk)
		if (`RST)	ready <= 0;
		else 		ready <= cnt_en;

	always @(posedge clk) begin
		if (cnt_en == 1'b0) begin
			dt	<=	1'b0;
		end
		else	begin	//1) W_1(66), 2) D_3(167), 3) N_13(166), 4) P_15(1666)
			case	(count)
				5'd0	:	begin
					case (cnt)
						10'd0	:	dt	<=	203	;
						10'd1	:	dt	<=	205	;
						10'd2	:	dt	<=	207	;
						10'd3	:	dt	<=	206	;
						10'd4	:	dt	<=	207	;
						10'd5	:	dt	<=	209	;
						10'd6	:	dt	<=	210	;
						10'd7	:	dt	<=	209	;
						10'd8	:	dt	<=	210	;
						10'd9	:	dt	<=	209	;
						10'd10	:	dt	<=	208	;
						10'd11	:	dt	<=	207	;
						10'd12	:	dt	<=	207	;
						10'd13	:	dt	<=	209	;
						10'd14	:	dt	<=	208	;
						10'd15	:	dt	<=	210	;
						10'd16	:	dt	<=	210	;
						10'd17	:	dt	<=	207	;
						10'd18	:	dt	<=	209	;
						10'd19	:	dt	<=	209	;
						10'd20	:	dt	<=	208	;
						10'd21	:	dt	<=	209	;
						10'd22	:	dt	<=	210	;
						10'd23	:	dt	<=	209	;
						10'd24	:	dt	<=	207	;
						10'd25	:	dt	<=	208	;
						10'd26	:	dt	<=	209	;
						10'd27	:	dt	<=	207	;
						10'd28	:	dt	<=	206	;
						10'd29	:	dt	<=	208	;
						10'd30	:	dt	<=	209	;
						10'd31	:	dt	<=	208	;
						10'd32	:	dt	<=	208	;
						10'd33	:	dt	<=	210	;
						10'd34	:	dt	<=	211	;
						10'd35	:	dt	<=	210	;
						10'd36	:	dt	<=	211	;
						10'd37	:	dt	<=	209	;
						10'd38	:	dt	<=	209	;
						10'd39	:	dt	<=	210	;
						10'd40	:	dt	<=	211	;
						10'd41	:	dt	<=	211	;
						10'd42	:	dt	<=	209	;
						10'd43	:	dt	<=	208	;
						10'd44	:	dt	<=	211	;
						10'd45	:	dt	<=	215	;
						10'd46	:	dt	<=	210	;
						10'd47	:	dt	<=	212	;
						10'd48	:	dt	<=	212	;
						10'd49	:	dt	<=	211	;
						10'd50	:	dt	<=	211	;
						10'd51	:	dt	<=	210	;
						10'd52	:	dt	<=	210	;
						10'd53	:	dt	<=	211	;
						10'd54	:	dt	<=	210	;
						10'd55	:	dt	<=	210	;
						10'd56	:	dt	<=	209	;
						10'd57	:	dt	<=	209	;
						10'd58	:	dt	<=	210	;
						10'd59	:	dt	<=	211	;
						10'd60	:	dt	<=	210	;
						10'd61	:	dt	<=	210	;
						10'd62	:	dt	<=	212	;
						10'd63	:	dt	<=	212	;
						10'd64	:	dt	<=	211	;
						10'd65	:	dt	<=	212	;
						10'd66	:	dt	<=	210	;
						10'd67	:	dt	<=	210	;
						10'd68	:	dt	<=	212	;
						10'd69	:	dt	<=	211	;
						10'd70	:	dt	<=	223	;
						10'd71	:	dt	<=	208	;
						10'd72	:	dt	<=	162	;
						10'd73	:	dt	<=	176	;
						10'd74	:	dt	<=	219	;
						10'd75	:	dt	<=	204	;
						10'd76	:	dt	<=	206	;
						10'd77	:	dt	<=	217	;
						10'd78	:	dt	<=	216	;
						10'd79	:	dt	<=	214	;
						10'd80	:	dt	<=	212	;
						10'd81	:	dt	<=	209	;
						10'd82	:	dt	<=	211	;
						10'd83	:	dt	<=	212	;
						10'd84	:	dt	<=	209	;
						10'd85	:	dt	<=	210	;
						10'd86	:	dt	<=	211	;
						10'd87	:	dt	<=	213	;
						10'd88	:	dt	<=	215	;
						10'd89	:	dt	<=	213	;
						10'd90	:	dt	<=	211	;
						10'd91	:	dt	<=	213	;
						10'd92	:	dt	<=	213	;
						10'd93	:	dt	<=	211	;
						10'd94	:	dt	<=	216	;
						10'd95	:	dt	<=	216	;
						10'd96	:	dt	<=	179	;
						10'd97	:	dt	<=	167	;
						10'd98	:	dt	<=	228	;
						10'd99	:	dt	<=	202	;
						10'd100	:	dt	<=	161	;
						10'd101	:	dt	<=	129	;
						10'd102	:	dt	<=	132	;
						10'd103	:	dt	<=	155	;
						10'd104	:	dt	<=	141	;
						10'd105	:	dt	<=	187	;
						10'd106	:	dt	<=	210	;
						10'd107	:	dt	<=	159	;
						10'd108	:	dt	<=	197	;
						10'd109	:	dt	<=	217	;
						10'd110	:	dt	<=	211	;
						10'd111	:	dt	<=	211	;
						10'd112	:	dt	<=	210	;
						10'd113	:	dt	<=	211	;
						10'd114	:	dt	<=	211	;
						10'd115	:	dt	<=	213	;
						10'd116	:	dt	<=	214	;
						10'd117	:	dt	<=	213	;
						10'd118	:	dt	<=	213	;
						10'd119	:	dt	<=	214	;
						10'd120	:	dt	<=	215	;
						10'd121	:	dt	<=	216	;
						10'd122	:	dt	<=	245	;
						10'd123	:	dt	<=	228	;
						10'd124	:	dt	<=	181	;
						10'd125	:	dt	<=	138	;
						10'd126	:	dt	<=	184	;
						10'd127	:	dt	<=	210	;
						10'd128	:	dt	<=	175	;
						10'd129	:	dt	<=	160	;
						10'd130	:	dt	<=	76	;
						10'd131	:	dt	<=	133	;
						10'd132	:	dt	<=	143	;
						10'd133	:	dt	<=	118	;
						10'd134	:	dt	<=	180	;
						10'd135	:	dt	<=	126	;
						10'd136	:	dt	<=	170	;
						10'd137	:	dt	<=	225	;
						10'd138	:	dt	<=	211	;
						10'd139	:	dt	<=	214	;
						10'd140	:	dt	<=	210	;
						10'd141	:	dt	<=	212	;
						10'd142	:	dt	<=	213	;
						10'd143	:	dt	<=	213	;
						10'd144	:	dt	<=	213	;
						10'd145	:	dt	<=	215	;
						10'd146	:	dt	<=	213	;
						10'd147	:	dt	<=	221	;
						10'd148	:	dt	<=	198	;
						10'd149	:	dt	<=	181	;
						10'd150	:	dt	<=	245	;
						10'd151	:	dt	<=	225	;
						10'd152	:	dt	<=	192	;
						10'd153	:	dt	<=	156	;
						10'd154	:	dt	<=	176	;
						10'd155	:	dt	<=	234	;
						10'd156	:	dt	<=	181	;
						10'd157	:	dt	<=	168	;
						10'd158	:	dt	<=	95	;
						10'd159	:	dt	<=	158	;
						10'd160	:	dt	<=	159	;
						10'd161	:	dt	<=	121	;
						10'd162	:	dt	<=	145	;
						10'd163	:	dt	<=	134	;
						10'd164	:	dt	<=	161	;
						10'd165	:	dt	<=	228	;
						10'd166	:	dt	<=	214	;
						10'd167	:	dt	<=	216	;
						10'd168	:	dt	<=	211	;
						10'd169	:	dt	<=	213	;
						10'd170	:	dt	<=	214	;
						10'd171	:	dt	<=	215	;
						10'd172	:	dt	<=	215	;
						10'd173	:	dt	<=	215	;
						10'd174	:	dt	<=	218	;
						10'd175	:	dt	<=	252	;
						10'd176	:	dt	<=	199	;
						10'd177	:	dt	<=	142	;
						10'd178	:	dt	<=	192	;
						10'd179	:	dt	<=	244	;
						10'd180	:	dt	<=	200	;
						10'd181	:	dt	<=	166	;
						10'd182	:	dt	<=	160	;
						10'd183	:	dt	<=	249	;
						10'd184	:	dt	<=	199	;
						10'd185	:	dt	<=	175	;
						10'd186	:	dt	<=	102	;
						10'd187	:	dt	<=	176	;
						10'd188	:	dt	<=	164	;
						10'd189	:	dt	<=	113	;
						10'd190	:	dt	<=	111	;
						10'd191	:	dt	<=	137	;
						10'd192	:	dt	<=	131	;
						10'd193	:	dt	<=	232	;
						10'd194	:	dt	<=	213	;
						10'd195	:	dt	<=	217	;
						10'd196	:	dt	<=	213	;
						10'd197	:	dt	<=	214	;
						10'd198	:	dt	<=	214	;
						10'd199	:	dt	<=	215	;
						10'd200	:	dt	<=	217	;
						10'd201	:	dt	<=	211	;
						10'd202	:	dt	<=	235	;
						10'd203	:	dt	<=	246	;
						10'd204	:	dt	<=	207	;
						10'd205	:	dt	<=	174	;
						10'd206	:	dt	<=	164	;
						10'd207	:	dt	<=	250	;
						10'd208	:	dt	<=	211	;
						10'd209	:	dt	<=	166	;
						10'd210	:	dt	<=	144	;
						10'd211	:	dt	<=	248	;
						10'd212	:	dt	<=	204	;
						10'd213	:	dt	<=	171	;
						10'd214	:	dt	<=	96	;
						10'd215	:	dt	<=	179	;
						10'd216	:	dt	<=	161	;
						10'd217	:	dt	<=	98	;
						10'd218	:	dt	<=	94	;
						10'd219	:	dt	<=	152	;
						10'd220	:	dt	<=	85	;
						10'd221	:	dt	<=	209	;
						10'd222	:	dt	<=	221	;
						10'd223	:	dt	<=	217	;
						10'd224	:	dt	<=	214	;
						10'd225	:	dt	<=	216	;
						10'd226	:	dt	<=	216	;
						10'd227	:	dt	<=	216	;
						10'd228	:	dt	<=	214	;
						10'd229	:	dt	<=	233	;
						10'd230	:	dt	<=	229	;
						10'd231	:	dt	<=	227	;
						10'd232	:	dt	<=	222	;
						10'd233	:	dt	<=	190	;
						10'd234	:	dt	<=	140	;
						10'd235	:	dt	<=	226	;
						10'd236	:	dt	<=	220	;
						10'd237	:	dt	<=	160	;
						10'd238	:	dt	<=	123	;
						10'd239	:	dt	<=	239	;
						10'd240	:	dt	<=	206	;
						10'd241	:	dt	<=	155	;
						10'd242	:	dt	<=	77	;
						10'd243	:	dt	<=	138	;
						10'd244	:	dt	<=	144	;
						10'd245	:	dt	<=	88	;
						10'd246	:	dt	<=	82	;
						10'd247	:	dt	<=	161	;
						10'd248	:	dt	<=	76	;
						10'd249	:	dt	<=	141	;
						10'd250	:	dt	<=	233	;
						10'd251	:	dt	<=	216	;
						10'd252	:	dt	<=	215	;
						10'd253	:	dt	<=	216	;
						10'd254	:	dt	<=	217	;
						10'd255	:	dt	<=	216	;
						10'd256	:	dt	<=	217	;
						10'd257	:	dt	<=	237	;
						10'd258	:	dt	<=	194	;
						10'd259	:	dt	<=	217	;
						10'd260	:	dt	<=	235	;
						10'd261	:	dt	<=	197	;
						10'd262	:	dt	<=	131	;
						10'd263	:	dt	<=	193	;
						10'd264	:	dt	<=	228	;
						10'd265	:	dt	<=	158	;
						10'd266	:	dt	<=	100	;
						10'd267	:	dt	<=	198	;
						10'd268	:	dt	<=	194	;
						10'd269	:	dt	<=	137	;
						10'd270	:	dt	<=	69	;
						10'd271	:	dt	<=	105	;
						10'd272	:	dt	<=	127	;
						10'd273	:	dt	<=	78	;
						10'd274	:	dt	<=	84	;
						10'd275	:	dt	<=	166	;
						10'd276	:	dt	<=	89	;
						10'd277	:	dt	<=	111	;
						10'd278	:	dt	<=	231	;
						10'd279	:	dt	<=	218	;
						10'd280	:	dt	<=	217	;
						10'd281	:	dt	<=	217	;
						10'd282	:	dt	<=	219	;
						10'd283	:	dt	<=	214	;
						10'd284	:	dt	<=	230	;
						10'd285	:	dt	<=	230	;
						10'd286	:	dt	<=	180	;
						10'd287	:	dt	<=	192	;
						10'd288	:	dt	<=	229	;
						10'd289	:	dt	<=	195	;
						10'd290	:	dt	<=	129	;
						10'd291	:	dt	<=	156	;
						10'd292	:	dt	<=	217	;
						10'd293	:	dt	<=	151	;
						10'd294	:	dt	<=	87	;
						10'd295	:	dt	<=	153	;
						10'd296	:	dt	<=	177	;
						10'd297	:	dt	<=	128	;
						10'd298	:	dt	<=	78	;
						10'd299	:	dt	<=	88	;
						10'd300	:	dt	<=	114	;
						10'd301	:	dt	<=	64	;
						10'd302	:	dt	<=	102	;
						10'd303	:	dt	<=	178	;
						10'd304	:	dt	<=	106	;
						10'd305	:	dt	<=	115	;
						10'd306	:	dt	<=	233	;
						10'd307	:	dt	<=	220	;
						10'd308	:	dt	<=	217	;
						10'd309	:	dt	<=	218	;
						10'd310	:	dt	<=	218	;
						10'd311	:	dt	<=	216	;
						10'd312	:	dt	<=	230	;
						10'd313	:	dt	<=	223	;
						10'd314	:	dt	<=	188	;
						10'd315	:	dt	<=	176	;
						10'd316	:	dt	<=	204	;
						10'd317	:	dt	<=	173	;
						10'd318	:	dt	<=	118	;
						10'd319	:	dt	<=	121	;
						10'd320	:	dt	<=	191	;
						10'd321	:	dt	<=	141	;
						10'd322	:	dt	<=	81	;
						10'd323	:	dt	<=	110	;
						10'd324	:	dt	<=	168	;
						10'd325	:	dt	<=	123	;
						10'd326	:	dt	<=	74	;
						10'd327	:	dt	<=	88	;
						10'd328	:	dt	<=	117	;
						10'd329	:	dt	<=	74	;
						10'd330	:	dt	<=	157	;
						10'd331	:	dt	<=	195	;
						10'd332	:	dt	<=	120	;
						10'd333	:	dt	<=	119	;
						10'd334	:	dt	<=	234	;
						10'd335	:	dt	<=	222	;
						10'd336	:	dt	<=	213	;
						10'd337	:	dt	<=	216	;
						10'd338	:	dt	<=	215	;
						10'd339	:	dt	<=	221	;
						10'd340	:	dt	<=	232	;
						10'd341	:	dt	<=	209	;
						10'd342	:	dt	<=	174	;
						10'd343	:	dt	<=	140	;
						10'd344	:	dt	<=	183	;
						10'd345	:	dt	<=	167	;
						10'd346	:	dt	<=	113	;
						10'd347	:	dt	<=	96	;
						10'd348	:	dt	<=	178	;
						10'd349	:	dt	<=	139	;
						10'd350	:	dt	<=	71	;
						10'd351	:	dt	<=	82	;
						10'd352	:	dt	<=	166	;
						10'd353	:	dt	<=	122	;
						10'd354	:	dt	<=	64	;
						10'd355	:	dt	<=	111	;
						10'd356	:	dt	<=	127	;
						10'd357	:	dt	<=	97	;
						10'd358	:	dt	<=	196	;
						10'd359	:	dt	<=	189	;
						10'd360	:	dt	<=	122	;
						10'd361	:	dt	<=	128	;
						10'd362	:	dt	<=	235	;
						10'd363	:	dt	<=	221	;
						10'd364	:	dt	<=	213	;
						10'd365	:	dt	<=	215	;
						10'd366	:	dt	<=	215	;
						10'd367	:	dt	<=	215	;
						10'd368	:	dt	<=	246	;
						10'd369	:	dt	<=	229	;
						10'd370	:	dt	<=	187	;
						10'd371	:	dt	<=	129	;
						10'd372	:	dt	<=	145	;
						10'd373	:	dt	<=	170	;
						10'd374	:	dt	<=	101	;
						10'd375	:	dt	<=	83	;
						10'd376	:	dt	<=	169	;
						10'd377	:	dt	<=	144	;
						10'd378	:	dt	<=	70	;
						10'd379	:	dt	<=	75	;
						10'd380	:	dt	<=	173	;
						10'd381	:	dt	<=	120	;
						10'd382	:	dt	<=	130	;
						10'd383	:	dt	<=	197	;
						10'd384	:	dt	<=	163	;
						10'd385	:	dt	<=	118	;
						10'd386	:	dt	<=	184	;
						10'd387	:	dt	<=	196	;
						10'd388	:	dt	<=	122	;
						10'd389	:	dt	<=	138	;
						10'd390	:	dt	<=	234	;
						10'd391	:	dt	<=	220	;
						10'd392	:	dt	<=	215	;
						10'd393	:	dt	<=	217	;
						10'd394	:	dt	<=	216	;
						10'd395	:	dt	<=	217	;
						10'd396	:	dt	<=	244	;
						10'd397	:	dt	<=	231	;
						10'd398	:	dt	<=	192	;
						10'd399	:	dt	<=	146	;
						10'd400	:	dt	<=	100	;
						10'd401	:	dt	<=	141	;
						10'd402	:	dt	<=	131	;
						10'd403	:	dt	<=	79	;
						10'd404	:	dt	<=	171	;
						10'd405	:	dt	<=	165	;
						10'd406	:	dt	<=	82	;
						10'd407	:	dt	<=	85	;
						10'd408	:	dt	<=	170	;
						10'd409	:	dt	<=	173	;
						10'd410	:	dt	<=	196	;
						10'd411	:	dt	<=	194	;
						10'd412	:	dt	<=	173	;
						10'd413	:	dt	<=	137	;
						10'd414	:	dt	<=	132	;
						10'd415	:	dt	<=	180	;
						10'd416	:	dt	<=	112	;
						10'd417	:	dt	<=	145	;
						10'd418	:	dt	<=	236	;
						10'd419	:	dt	<=	221	;
						10'd420	:	dt	<=	217	;
						10'd421	:	dt	<=	218	;
						10'd422	:	dt	<=	217	;
						10'd423	:	dt	<=	221	;
						10'd424	:	dt	<=	248	;
						10'd425	:	dt	<=	235	;
						10'd426	:	dt	<=	206	;
						10'd427	:	dt	<=	169	;
						10'd428	:	dt	<=	123	;
						10'd429	:	dt	<=	109	;
						10'd430	:	dt	<=	140	;
						10'd431	:	dt	<=	103	;
						10'd432	:	dt	<=	164	;
						10'd433	:	dt	<=	178	;
						10'd434	:	dt	<=	148	;
						10'd435	:	dt	<=	189	;
						10'd436	:	dt	<=	206	;
						10'd437	:	dt	<=	203	;
						10'd438	:	dt	<=	191	;
						10'd439	:	dt	<=	177	;
						10'd440	:	dt	<=	154	;
						10'd441	:	dt	<=	137	;
						10'd442	:	dt	<=	114	;
						10'd443	:	dt	<=	117	;
						10'd444	:	dt	<=	91	;
						10'd445	:	dt	<=	138	;
						10'd446	:	dt	<=	238	;
						10'd447	:	dt	<=	220	;
						10'd448	:	dt	<=	218	;
						10'd449	:	dt	<=	219	;
						10'd450	:	dt	<=	219	;
						10'd451	:	dt	<=	221	;
						10'd452	:	dt	<=	249	;
						10'd453	:	dt	<=	243	;
						10'd454	:	dt	<=	214	;
						10'd455	:	dt	<=	182	;
						10'd456	:	dt	<=	164	;
						10'd457	:	dt	<=	151	;
						10'd458	:	dt	<=	142	;
						10'd459	:	dt	<=	164	;
						10'd460	:	dt	<=	185	;
						10'd461	:	dt	<=	198	;
						10'd462	:	dt	<=	218	;
						10'd463	:	dt	<=	220	;
						10'd464	:	dt	<=	218	;
						10'd465	:	dt	<=	207	;
						10'd466	:	dt	<=	189	;
						10'd467	:	dt	<=	170	;
						10'd468	:	dt	<=	143	;
						10'd469	:	dt	<=	121	;
						10'd470	:	dt	<=	113	;
						10'd471	:	dt	<=	92	;
						10'd472	:	dt	<=	73	;
						10'd473	:	dt	<=	131	;
						10'd474	:	dt	<=	239	;
						10'd475	:	dt	<=	220	;
						10'd476	:	dt	<=	217	;
						10'd477	:	dt	<=	218	;
						10'd478	:	dt	<=	217	;
						10'd479	:	dt	<=	222	;
						10'd480	:	dt	<=	244	;
						10'd481	:	dt	<=	243	;
						10'd482	:	dt	<=	223	;
						10'd483	:	dt	<=	200	;
						10'd484	:	dt	<=	185	;
						10'd485	:	dt	<=	173	;
						10'd486	:	dt	<=	160	;
						10'd487	:	dt	<=	160	;
						10'd488	:	dt	<=	187	;
						10'd489	:	dt	<=	205	;
						10'd490	:	dt	<=	218	;
						10'd491	:	dt	<=	217	;
						10'd492	:	dt	<=	218	;
						10'd493	:	dt	<=	209	;
						10'd494	:	dt	<=	183	;
						10'd495	:	dt	<=	164	;
						10'd496	:	dt	<=	142	;
						10'd497	:	dt	<=	114	;
						10'd498	:	dt	<=	99	;
						10'd499	:	dt	<=	93	;
						10'd500	:	dt	<=	66	;
						10'd501	:	dt	<=	159	;
						10'd502	:	dt	<=	238	;
						10'd503	:	dt	<=	222	;
						10'd504	:	dt	<=	216	;
						10'd505	:	dt	<=	216	;
						10'd506	:	dt	<=	217	;
						10'd507	:	dt	<=	221	;
						10'd508	:	dt	<=	238	;
						10'd509	:	dt	<=	238	;
						10'd510	:	dt	<=	231	;
						10'd511	:	dt	<=	215	;
						10'd512	:	dt	<=	204	;
						10'd513	:	dt	<=	182	;
						10'd514	:	dt	<=	170	;
						10'd515	:	dt	<=	165	;
						10'd516	:	dt	<=	178	;
						10'd517	:	dt	<=	201	;
						10'd518	:	dt	<=	215	;
						10'd519	:	dt	<=	216	;
						10'd520	:	dt	<=	211	;
						10'd521	:	dt	<=	202	;
						10'd522	:	dt	<=	177	;
						10'd523	:	dt	<=	157	;
						10'd524	:	dt	<=	136	;
						10'd525	:	dt	<=	110	;
						10'd526	:	dt	<=	96	;
						10'd527	:	dt	<=	76	;
						10'd528	:	dt	<=	113	;
						10'd529	:	dt	<=	222	;
						10'd530	:	dt	<=	230	;
						10'd531	:	dt	<=	227	;
						10'd532	:	dt	<=	222	;
						10'd533	:	dt	<=	223	;
						10'd534	:	dt	<=	224	;
						10'd535	:	dt	<=	216	;
						10'd536	:	dt	<=	233	;
						10'd537	:	dt	<=	239	;
						10'd538	:	dt	<=	240	;
						10'd539	:	dt	<=	229	;
						10'd540	:	dt	<=	210	;
						10'd541	:	dt	<=	187	;
						10'd542	:	dt	<=	171	;
						10'd543	:	dt	<=	168	;
						10'd544	:	dt	<=	180	;
						10'd545	:	dt	<=	207	;
						10'd546	:	dt	<=	218	;
						10'd547	:	dt	<=	218	;
						10'd548	:	dt	<=	203	;
						10'd549	:	dt	<=	194	;
						10'd550	:	dt	<=	174	;
						10'd551	:	dt	<=	153	;
						10'd552	:	dt	<=	129	;
						10'd553	:	dt	<=	107	;
						10'd554	:	dt	<=	80	;
						10'd555	:	dt	<=	97	;
						10'd556	:	dt	<=	213	;
						10'd557	:	dt	<=	227	;
						10'd558	:	dt	<=	225	;
						10'd559	:	dt	<=	226	;
						10'd560	:	dt	<=	175	;
						10'd561	:	dt	<=	180	;
						10'd562	:	dt	<=	188	;
						10'd563	:	dt	<=	178	;
						10'd564	:	dt	<=	214	;
						10'd565	:	dt	<=	240	;
						10'd566	:	dt	<=	245	;
						10'd567	:	dt	<=	233	;
						10'd568	:	dt	<=	210	;
						10'd569	:	dt	<=	191	;
						10'd570	:	dt	<=	174	;
						10'd571	:	dt	<=	167	;
						10'd572	:	dt	<=	179	;
						10'd573	:	dt	<=	211	;
						10'd574	:	dt	<=	220	;
						10'd575	:	dt	<=	211	;
						10'd576	:	dt	<=	196	;
						10'd577	:	dt	<=	186	;
						10'd578	:	dt	<=	168	;
						10'd579	:	dt	<=	143	;
						10'd580	:	dt	<=	118	;
						10'd581	:	dt	<=	96	;
						10'd582	:	dt	<=	78	;
						10'd583	:	dt	<=	196	;
						10'd584	:	dt	<=	239	;
						10'd585	:	dt	<=	230	;
						10'd586	:	dt	<=	234	;
						10'd587	:	dt	<=	233	;
						10'd588	:	dt	<=	94	;
						10'd589	:	dt	<=	96	;
						10'd590	:	dt	<=	103	;
						10'd591	:	dt	<=	85	;
						10'd592	:	dt	<=	151	;
						10'd593	:	dt	<=	244	;
						10'd594	:	dt	<=	234	;
						10'd595	:	dt	<=	226	;
						10'd596	:	dt	<=	211	;
						10'd597	:	dt	<=	195	;
						10'd598	:	dt	<=	181	;
						10'd599	:	dt	<=	165	;
						10'd600	:	dt	<=	178	;
						10'd601	:	dt	<=	207	;
						10'd602	:	dt	<=	207	;
						10'd603	:	dt	<=	192	;
						10'd604	:	dt	<=	178	;
						10'd605	:	dt	<=	168	;
						10'd606	:	dt	<=	153	;
						10'd607	:	dt	<=	129	;
						10'd608	:	dt	<=	107	;
						10'd609	:	dt	<=	86	;
						10'd610	:	dt	<=	104	;
						10'd611	:	dt	<=	177	;
						10'd612	:	dt	<=	178	;
						10'd613	:	dt	<=	182	;
						10'd614	:	dt	<=	178	;
						10'd615	:	dt	<=	177	;
						10'd616	:	dt	<=	103	;
						10'd617	:	dt	<=	103	;
						10'd618	:	dt	<=	104	;
						10'd619	:	dt	<=	91	;
						10'd620	:	dt	<=	114	;
						10'd621	:	dt	<=	239	;
						10'd622	:	dt	<=	220	;
						10'd623	:	dt	<=	212	;
						10'd624	:	dt	<=	211	;
						10'd625	:	dt	<=	202	;
						10'd626	:	dt	<=	188	;
						10'd627	:	dt	<=	164	;
						10'd628	:	dt	<=	173	;
						10'd629	:	dt	<=	203	;
						10'd630	:	dt	<=	198	;
						10'd631	:	dt	<=	178	;
						10'd632	:	dt	<=	156	;
						10'd633	:	dt	<=	140	;
						10'd634	:	dt	<=	127	;
						10'd635	:	dt	<=	115	;
						10'd636	:	dt	<=	95	;
						10'd637	:	dt	<=	92	;
						10'd638	:	dt	<=	99	;
						10'd639	:	dt	<=	95	;
						10'd640	:	dt	<=	90	;
						10'd641	:	dt	<=	86	;
						10'd642	:	dt	<=	113	;
						10'd643	:	dt	<=	156	;
						10'd644	:	dt	<=	101	;
						10'd645	:	dt	<=	103	;
						10'd646	:	dt	<=	105	;
						10'd647	:	dt	<=	99	;
						10'd648	:	dt	<=	106	;
						10'd649	:	dt	<=	230	;
						10'd650	:	dt	<=	209	;
						10'd651	:	dt	<=	204	;
						10'd652	:	dt	<=	214	;
						10'd653	:	dt	<=	204	;
						10'd654	:	dt	<=	185	;
						10'd655	:	dt	<=	164	;
						10'd656	:	dt	<=	167	;
						10'd657	:	dt	<=	201	;
						10'd658	:	dt	<=	194	;
						10'd659	:	dt	<=	168	;
						10'd660	:	dt	<=	131	;
						10'd661	:	dt	<=	109	;
						10'd662	:	dt	<=	103	;
						10'd663	:	dt	<=	93	;
						10'd664	:	dt	<=	93	;
						10'd665	:	dt	<=	104	;
						10'd666	:	dt	<=	98	;
						10'd667	:	dt	<=	97	;
						10'd668	:	dt	<=	131	;
						10'd669	:	dt	<=	187	;
						10'd670	:	dt	<=	234	;
						10'd671	:	dt	<=	233	;
						10'd672	:	dt	<=	100	;
						10'd673	:	dt	<=	101	;
						10'd674	:	dt	<=	100	;
						10'd675	:	dt	<=	102	;
						10'd676	:	dt	<=	104	;
						10'd677	:	dt	<=	222	;
						10'd678	:	dt	<=	207	;
						10'd679	:	dt	<=	205	;
						10'd680	:	dt	<=	215	;
						10'd681	:	dt	<=	199	;
						10'd682	:	dt	<=	183	;
						10'd683	:	dt	<=	172	;
						10'd684	:	dt	<=	164	;
						10'd685	:	dt	<=	193	;
						10'd686	:	dt	<=	187	;
						10'd687	:	dt	<=	153	;
						10'd688	:	dt	<=	107	;
						10'd689	:	dt	<=	91	;
						10'd690	:	dt	<=	86	;
						10'd691	:	dt	<=	93	;
						10'd692	:	dt	<=	102	;
						10'd693	:	dt	<=	108	;
						10'd694	:	dt	<=	141	;
						10'd695	:	dt	<=	195	;
						10'd696	:	dt	<=	241	;
						10'd697	:	dt	<=	242	;
						10'd698	:	dt	<=	226	;
						10'd699	:	dt	<=	207	;
						10'd700	:	dt	<=	100	;
						10'd701	:	dt	<=	101	;
						10'd702	:	dt	<=	100	;
						10'd703	:	dt	<=	104	;
					endcase
				end
				5'd1	:	begin
					case (cnt)
						10'd0	:	dt	<=	92	;
						10'd1	:	dt	<=	95	;
						10'd2	:	dt	<=	82	;
						10'd3	:	dt	<=	69	;
						10'd4	:	dt	<=	65	;
						10'd5	:	dt	<=	61	;
						10'd6	:	dt	<=	60	;
						10'd7	:	dt	<=	34	;
						10'd8	:	dt	<=	54	;
						10'd9	:	dt	<=	81	;
						10'd10	:	dt	<=	97	;
						10'd11	:	dt	<=	112	;
						10'd12	:	dt	<=	135	;
						10'd13	:	dt	<=	118	;
						10'd14	:	dt	<=	105	;
						10'd15	:	dt	<=	125	;
						10'd16	:	dt	<=	129	;
						10'd17	:	dt	<=	136	;
						10'd18	:	dt	<=	141	;
						10'd19	:	dt	<=	144	;
						10'd20	:	dt	<=	147	;
						10'd21	:	dt	<=	150	;
						10'd22	:	dt	<=	152	;
						10'd23	:	dt	<=	154	;
						10'd24	:	dt	<=	156	;
						10'd25	:	dt	<=	157	;
						10'd26	:	dt	<=	159	;
						10'd27	:	dt	<=	160	;
						10'd28	:	dt	<=	94	;
						10'd29	:	dt	<=	97	;
						10'd30	:	dt	<=	82	;
						10'd31	:	dt	<=	70	;
						10'd32	:	dt	<=	65	;
						10'd33	:	dt	<=	64	;
						10'd34	:	dt	<=	60	;
						10'd35	:	dt	<=	35	;
						10'd36	:	dt	<=	58	;
						10'd37	:	dt	<=	84	;
						10'd38	:	dt	<=	104	;
						10'd39	:	dt	<=	116	;
						10'd40	:	dt	<=	136	;
						10'd41	:	dt	<=	124	;
						10'd42	:	dt	<=	102	;
						10'd43	:	dt	<=	122	;
						10'd44	:	dt	<=	115	;
						10'd45	:	dt	<=	126	;
						10'd46	:	dt	<=	142	;
						10'd47	:	dt	<=	145	;
						10'd48	:	dt	<=	148	;
						10'd49	:	dt	<=	151	;
						10'd50	:	dt	<=	153	;
						10'd51	:	dt	<=	156	;
						10'd52	:	dt	<=	157	;
						10'd53	:	dt	<=	158	;
						10'd54	:	dt	<=	160	;
						10'd55	:	dt	<=	161	;
						10'd56	:	dt	<=	97	;
						10'd57	:	dt	<=	98	;
						10'd58	:	dt	<=	81	;
						10'd59	:	dt	<=	72	;
						10'd60	:	dt	<=	65	;
						10'd61	:	dt	<=	67	;
						10'd62	:	dt	<=	57	;
						10'd63	:	dt	<=	36	;
						10'd64	:	dt	<=	62	;
						10'd65	:	dt	<=	88	;
						10'd66	:	dt	<=	122	;
						10'd67	:	dt	<=	122	;
						10'd68	:	dt	<=	126	;
						10'd69	:	dt	<=	132	;
						10'd70	:	dt	<=	109	;
						10'd71	:	dt	<=	129	;
						10'd72	:	dt	<=	112	;
						10'd73	:	dt	<=	111	;
						10'd74	:	dt	<=	140	;
						10'd75	:	dt	<=	147	;
						10'd76	:	dt	<=	150	;
						10'd77	:	dt	<=	152	;
						10'd78	:	dt	<=	154	;
						10'd79	:	dt	<=	157	;
						10'd80	:	dt	<=	158	;
						10'd81	:	dt	<=	159	;
						10'd82	:	dt	<=	161	;
						10'd83	:	dt	<=	162	;
						10'd84	:	dt	<=	99	;
						10'd85	:	dt	<=	98	;
						10'd86	:	dt	<=	80	;
						10'd87	:	dt	<=	74	;
						10'd88	:	dt	<=	67	;
						10'd89	:	dt	<=	70	;
						10'd90	:	dt	<=	53	;
						10'd91	:	dt	<=	38	;
						10'd92	:	dt	<=	66	;
						10'd93	:	dt	<=	92	;
						10'd94	:	dt	<=	133	;
						10'd95	:	dt	<=	128	;
						10'd96	:	dt	<=	120	;
						10'd97	:	dt	<=	137	;
						10'd98	:	dt	<=	117	;
						10'd99	:	dt	<=	134	;
						10'd100	:	dt	<=	122	;
						10'd101	:	dt	<=	104	;
						10'd102	:	dt	<=	136	;
						10'd103	:	dt	<=	148	;
						10'd104	:	dt	<=	151	;
						10'd105	:	dt	<=	153	;
						10'd106	:	dt	<=	156	;
						10'd107	:	dt	<=	158	;
						10'd108	:	dt	<=	159	;
						10'd109	:	dt	<=	161	;
						10'd110	:	dt	<=	162	;
						10'd111	:	dt	<=	163	;
						10'd112	:	dt	<=	102	;
						10'd113	:	dt	<=	97	;
						10'd114	:	dt	<=	80	;
						10'd115	:	dt	<=	76	;
						10'd116	:	dt	<=	68	;
						10'd117	:	dt	<=	72	;
						10'd118	:	dt	<=	49	;
						10'd119	:	dt	<=	41	;
						10'd120	:	dt	<=	71	;
						10'd121	:	dt	<=	95	;
						10'd122	:	dt	<=	137	;
						10'd123	:	dt	<=	133	;
						10'd124	:	dt	<=	122	;
						10'd125	:	dt	<=	148	;
						10'd126	:	dt	<=	129	;
						10'd127	:	dt	<=	133	;
						10'd128	:	dt	<=	131	;
						10'd129	:	dt	<=	105	;
						10'd130	:	dt	<=	131	;
						10'd131	:	dt	<=	150	;
						10'd132	:	dt	<=	152	;
						10'd133	:	dt	<=	155	;
						10'd134	:	dt	<=	157	;
						10'd135	:	dt	<=	159	;
						10'd136	:	dt	<=	161	;
						10'd137	:	dt	<=	163	;
						10'd138	:	dt	<=	164	;
						10'd139	:	dt	<=	165	;
						10'd140	:	dt	<=	104	;
						10'd141	:	dt	<=	97	;
						10'd142	:	dt	<=	81	;
						10'd143	:	dt	<=	78	;
						10'd144	:	dt	<=	70	;
						10'd145	:	dt	<=	74	;
						10'd146	:	dt	<=	46	;
						10'd147	:	dt	<=	45	;
						10'd148	:	dt	<=	77	;
						10'd149	:	dt	<=	99	;
						10'd150	:	dt	<=	138	;
						10'd151	:	dt	<=	139	;
						10'd152	:	dt	<=	126	;
						10'd153	:	dt	<=	155	;
						10'd154	:	dt	<=	136	;
						10'd155	:	dt	<=	134	;
						10'd156	:	dt	<=	145	;
						10'd157	:	dt	<=	113	;
						10'd158	:	dt	<=	125	;
						10'd159	:	dt	<=	151	;
						10'd160	:	dt	<=	155	;
						10'd161	:	dt	<=	157	;
						10'd162	:	dt	<=	159	;
						10'd163	:	dt	<=	161	;
						10'd164	:	dt	<=	163	;
						10'd165	:	dt	<=	165	;
						10'd166	:	dt	<=	166	;
						10'd167	:	dt	<=	167	;
						10'd168	:	dt	<=	107	;
						10'd169	:	dt	<=	97	;
						10'd170	:	dt	<=	84	;
						10'd171	:	dt	<=	81	;
						10'd172	:	dt	<=	72	;
						10'd173	:	dt	<=	76	;
						10'd174	:	dt	<=	43	;
						10'd175	:	dt	<=	51	;
						10'd176	:	dt	<=	98	;
						10'd177	:	dt	<=	113	;
						10'd178	:	dt	<=	139	;
						10'd179	:	dt	<=	149	;
						10'd180	:	dt	<=	129	;
						10'd181	:	dt	<=	152	;
						10'd182	:	dt	<=	138	;
						10'd183	:	dt	<=	136	;
						10'd184	:	dt	<=	155	;
						10'd185	:	dt	<=	123	;
						10'd186	:	dt	<=	118	;
						10'd187	:	dt	<=	150	;
						10'd188	:	dt	<=	157	;
						10'd189	:	dt	<=	159	;
						10'd190	:	dt	<=	161	;
						10'd191	:	dt	<=	164	;
						10'd192	:	dt	<=	166	;
						10'd193	:	dt	<=	168	;
						10'd194	:	dt	<=	168	;
						10'd195	:	dt	<=	168	;
						10'd196	:	dt	<=	109	;
						10'd197	:	dt	<=	97	;
						10'd198	:	dt	<=	86	;
						10'd199	:	dt	<=	82	;
						10'd200	:	dt	<=	74	;
						10'd201	:	dt	<=	76	;
						10'd202	:	dt	<=	41	;
						10'd203	:	dt	<=	60	;
						10'd204	:	dt	<=	120	;
						10'd205	:	dt	<=	122	;
						10'd206	:	dt	<=	136	;
						10'd207	:	dt	<=	151	;
						10'd208	:	dt	<=	128	;
						10'd209	:	dt	<=	146	;
						10'd210	:	dt	<=	140	;
						10'd211	:	dt	<=	133	;
						10'd212	:	dt	<=	154	;
						10'd213	:	dt	<=	129	;
						10'd214	:	dt	<=	114	;
						10'd215	:	dt	<=	148	;
						10'd216	:	dt	<=	158	;
						10'd217	:	dt	<=	160	;
						10'd218	:	dt	<=	163	;
						10'd219	:	dt	<=	166	;
						10'd220	:	dt	<=	168	;
						10'd221	:	dt	<=	169	;
						10'd222	:	dt	<=	169	;
						10'd223	:	dt	<=	170	;
						10'd224	:	dt	<=	110	;
						10'd225	:	dt	<=	97	;
						10'd226	:	dt	<=	88	;
						10'd227	:	dt	<=	82	;
						10'd228	:	dt	<=	77	;
						10'd229	:	dt	<=	75	;
						10'd230	:	dt	<=	40	;
						10'd231	:	dt	<=	66	;
						10'd232	:	dt	<=	127	;
						10'd233	:	dt	<=	122	;
						10'd234	:	dt	<=	133	;
						10'd235	:	dt	<=	150	;
						10'd236	:	dt	<=	126	;
						10'd237	:	dt	<=	145	;
						10'd238	:	dt	<=	146	;
						10'd239	:	dt	<=	130	;
						10'd240	:	dt	<=	153	;
						10'd241	:	dt	<=	135	;
						10'd242	:	dt	<=	113	;
						10'd243	:	dt	<=	147	;
						10'd244	:	dt	<=	160	;
						10'd245	:	dt	<=	162	;
						10'd246	:	dt	<=	165	;
						10'd247	:	dt	<=	168	;
						10'd248	:	dt	<=	169	;
						10'd249	:	dt	<=	171	;
						10'd250	:	dt	<=	171	;
						10'd251	:	dt	<=	172	;
						10'd252	:	dt	<=	111	;
						10'd253	:	dt	<=	96	;
						10'd254	:	dt	<=	90	;
						10'd255	:	dt	<=	82	;
						10'd256	:	dt	<=	80	;
						10'd257	:	dt	<=	73	;
						10'd258	:	dt	<=	39	;
						10'd259	:	dt	<=	71	;
						10'd260	:	dt	<=	132	;
						10'd261	:	dt	<=	125	;
						10'd262	:	dt	<=	131	;
						10'd263	:	dt	<=	153	;
						10'd264	:	dt	<=	126	;
						10'd265	:	dt	<=	142	;
						10'd266	:	dt	<=	151	;
						10'd267	:	dt	<=	129	;
						10'd268	:	dt	<=	154	;
						10'd269	:	dt	<=	141	;
						10'd270	:	dt	<=	114	;
						10'd271	:	dt	<=	144	;
						10'd272	:	dt	<=	161	;
						10'd273	:	dt	<=	164	;
						10'd274	:	dt	<=	167	;
						10'd275	:	dt	<=	169	;
						10'd276	:	dt	<=	171	;
						10'd277	:	dt	<=	172	;
						10'd278	:	dt	<=	173	;
						10'd279	:	dt	<=	173	;
						10'd280	:	dt	<=	111	;
						10'd281	:	dt	<=	96	;
						10'd282	:	dt	<=	92	;
						10'd283	:	dt	<=	82	;
						10'd284	:	dt	<=	83	;
						10'd285	:	dt	<=	69	;
						10'd286	:	dt	<=	39	;
						10'd287	:	dt	<=	74	;
						10'd288	:	dt	<=	138	;
						10'd289	:	dt	<=	135	;
						10'd290	:	dt	<=	130	;
						10'd291	:	dt	<=	156	;
						10'd292	:	dt	<=	128	;
						10'd293	:	dt	<=	129	;
						10'd294	:	dt	<=	147	;
						10'd295	:	dt	<=	124	;
						10'd296	:	dt	<=	148	;
						10'd297	:	dt	<=	142	;
						10'd298	:	dt	<=	112	;
						10'd299	:	dt	<=	140	;
						10'd300	:	dt	<=	163	;
						10'd301	:	dt	<=	166	;
						10'd302	:	dt	<=	168	;
						10'd303	:	dt	<=	170	;
						10'd304	:	dt	<=	172	;
						10'd305	:	dt	<=	174	;
						10'd306	:	dt	<=	174	;
						10'd307	:	dt	<=	174	;
						10'd308	:	dt	<=	109	;
						10'd309	:	dt	<=	97	;
						10'd310	:	dt	<=	94	;
						10'd311	:	dt	<=	83	;
						10'd312	:	dt	<=	87	;
						10'd313	:	dt	<=	65	;
						10'd314	:	dt	<=	41	;
						10'd315	:	dt	<=	76	;
						10'd316	:	dt	<=	137	;
						10'd317	:	dt	<=	137	;
						10'd318	:	dt	<=	123	;
						10'd319	:	dt	<=	153	;
						10'd320	:	dt	<=	130	;
						10'd321	:	dt	<=	117	;
						10'd322	:	dt	<=	140	;
						10'd323	:	dt	<=	121	;
						10'd324	:	dt	<=	140	;
						10'd325	:	dt	<=	142	;
						10'd326	:	dt	<=	110	;
						10'd327	:	dt	<=	134	;
						10'd328	:	dt	<=	163	;
						10'd329	:	dt	<=	167	;
						10'd330	:	dt	<=	169	;
						10'd331	:	dt	<=	172	;
						10'd332	:	dt	<=	174	;
						10'd333	:	dt	<=	175	;
						10'd334	:	dt	<=	175	;
						10'd335	:	dt	<=	175	;
						10'd336	:	dt	<=	108	;
						10'd337	:	dt	<=	97	;
						10'd338	:	dt	<=	95	;
						10'd339	:	dt	<=	82	;
						10'd340	:	dt	<=	89	;
						10'd341	:	dt	<=	60	;
						10'd342	:	dt	<=	43	;
						10'd343	:	dt	<=	77	;
						10'd344	:	dt	<=	132	;
						10'd345	:	dt	<=	139	;
						10'd346	:	dt	<=	117	;
						10'd347	:	dt	<=	145	;
						10'd348	:	dt	<=	137	;
						10'd349	:	dt	<=	128	;
						10'd350	:	dt	<=	138	;
						10'd351	:	dt	<=	138	;
						10'd352	:	dt	<=	145	;
						10'd353	:	dt	<=	129	;
						10'd354	:	dt	<=	101	;
						10'd355	:	dt	<=	123	;
						10'd356	:	dt	<=	162	;
						10'd357	:	dt	<=	168	;
						10'd358	:	dt	<=	170	;
						10'd359	:	dt	<=	173	;
						10'd360	:	dt	<=	175	;
						10'd361	:	dt	<=	176	;
						10'd362	:	dt	<=	176	;
						10'd363	:	dt	<=	176	;
						10'd364	:	dt	<=	107	;
						10'd365	:	dt	<=	98	;
						10'd366	:	dt	<=	95	;
						10'd367	:	dt	<=	83	;
						10'd368	:	dt	<=	90	;
						10'd369	:	dt	<=	55	;
						10'd370	:	dt	<=	45	;
						10'd371	:	dt	<=	78	;
						10'd372	:	dt	<=	132	;
						10'd373	:	dt	<=	146	;
						10'd374	:	dt	<=	119	;
						10'd375	:	dt	<=	138	;
						10'd376	:	dt	<=	147	;
						10'd377	:	dt	<=	137	;
						10'd378	:	dt	<=	133	;
						10'd379	:	dt	<=	148	;
						10'd380	:	dt	<=	146	;
						10'd381	:	dt	<=	111	;
						10'd382	:	dt	<=	87	;
						10'd383	:	dt	<=	111	;
						10'd384	:	dt	<=	160	;
						10'd385	:	dt	<=	170	;
						10'd386	:	dt	<=	172	;
						10'd387	:	dt	<=	174	;
						10'd388	:	dt	<=	175	;
						10'd389	:	dt	<=	177	;
						10'd390	:	dt	<=	178	;
						10'd391	:	dt	<=	179	;
						10'd392	:	dt	<=	106	;
						10'd393	:	dt	<=	100	;
						10'd394	:	dt	<=	95	;
						10'd395	:	dt	<=	83	;
						10'd396	:	dt	<=	90	;
						10'd397	:	dt	<=	51	;
						10'd398	:	dt	<=	49	;
						10'd399	:	dt	<=	81	;
						10'd400	:	dt	<=	132	;
						10'd401	:	dt	<=	147	;
						10'd402	:	dt	<=	132	;
						10'd403	:	dt	<=	143	;
						10'd404	:	dt	<=	147	;
						10'd405	:	dt	<=	144	;
						10'd406	:	dt	<=	144	;
						10'd407	:	dt	<=	162	;
						10'd408	:	dt	<=	154	;
						10'd409	:	dt	<=	114	;
						10'd410	:	dt	<=	83	;
						10'd411	:	dt	<=	97	;
						10'd412	:	dt	<=	153	;
						10'd413	:	dt	<=	170	;
						10'd414	:	dt	<=	173	;
						10'd415	:	dt	<=	175	;
						10'd416	:	dt	<=	176	;
						10'd417	:	dt	<=	177	;
						10'd418	:	dt	<=	179	;
						10'd419	:	dt	<=	180	;
						10'd420	:	dt	<=	106	;
						10'd421	:	dt	<=	101	;
						10'd422	:	dt	<=	95	;
						10'd423	:	dt	<=	83	;
						10'd424	:	dt	<=	89	;
						10'd425	:	dt	<=	46	;
						10'd426	:	dt	<=	51	;
						10'd427	:	dt	<=	83	;
						10'd428	:	dt	<=	136	;
						10'd429	:	dt	<=	155	;
						10'd430	:	dt	<=	149	;
						10'd431	:	dt	<=	140	;
						10'd432	:	dt	<=	139	;
						10'd433	:	dt	<=	142	;
						10'd434	:	dt	<=	148	;
						10'd435	:	dt	<=	158	;
						10'd436	:	dt	<=	155	;
						10'd437	:	dt	<=	130	;
						10'd438	:	dt	<=	94	;
						10'd439	:	dt	<=	87	;
						10'd440	:	dt	<=	144	;
						10'd441	:	dt	<=	171	;
						10'd442	:	dt	<=	174	;
						10'd443	:	dt	<=	176	;
						10'd444	:	dt	<=	177	;
						10'd445	:	dt	<=	178	;
						10'd446	:	dt	<=	179	;
						10'd447	:	dt	<=	181	;
						10'd448	:	dt	<=	105	;
						10'd449	:	dt	<=	103	;
						10'd450	:	dt	<=	95	;
						10'd451	:	dt	<=	86	;
						10'd452	:	dt	<=	89	;
						10'd453	:	dt	<=	43	;
						10'd454	:	dt	<=	54	;
						10'd455	:	dt	<=	87	;
						10'd456	:	dt	<=	145	;
						10'd457	:	dt	<=	164	;
						10'd458	:	dt	<=	148	;
						10'd459	:	dt	<=	131	;
						10'd460	:	dt	<=	128	;
						10'd461	:	dt	<=	134	;
						10'd462	:	dt	<=	140	;
						10'd463	:	dt	<=	146	;
						10'd464	:	dt	<=	155	;
						10'd465	:	dt	<=	151	;
						10'd466	:	dt	<=	118	;
						10'd467	:	dt	<=	90	;
						10'd468	:	dt	<=	133	;
						10'd469	:	dt	<=	170	;
						10'd470	:	dt	<=	174	;
						10'd471	:	dt	<=	176	;
						10'd472	:	dt	<=	177	;
						10'd473	:	dt	<=	178	;
						10'd474	:	dt	<=	180	;
						10'd475	:	dt	<=	181	;
						10'd476	:	dt	<=	104	;
						10'd477	:	dt	<=	105	;
						10'd478	:	dt	<=	96	;
						10'd479	:	dt	<=	90	;
						10'd480	:	dt	<=	87	;
						10'd481	:	dt	<=	40	;
						10'd482	:	dt	<=	56	;
						10'd483	:	dt	<=	90	;
						10'd484	:	dt	<=	149	;
						10'd485	:	dt	<=	162	;
						10'd486	:	dt	<=	139	;
						10'd487	:	dt	<=	123	;
						10'd488	:	dt	<=	126	;
						10'd489	:	dt	<=	135	;
						10'd490	:	dt	<=	148	;
						10'd491	:	dt	<=	161	;
						10'd492	:	dt	<=	167	;
						10'd493	:	dt	<=	167	;
						10'd494	:	dt	<=	142	;
						10'd495	:	dt	<=	104	;
						10'd496	:	dt	<=	121	;
						10'd497	:	dt	<=	167	;
						10'd498	:	dt	<=	175	;
						10'd499	:	dt	<=	177	;
						10'd500	:	dt	<=	178	;
						10'd501	:	dt	<=	179	;
						10'd502	:	dt	<=	180	;
						10'd503	:	dt	<=	181	;
						10'd504	:	dt	<=	104	;
						10'd505	:	dt	<=	107	;
						10'd506	:	dt	<=	95	;
						10'd507	:	dt	<=	93	;
						10'd508	:	dt	<=	84	;
						10'd509	:	dt	<=	39	;
						10'd510	:	dt	<=	59	;
						10'd511	:	dt	<=	89	;
						10'd512	:	dt	<=	143	;
						10'd513	:	dt	<=	159	;
						10'd514	:	dt	<=	135	;
						10'd515	:	dt	<=	120	;
						10'd516	:	dt	<=	128	;
						10'd517	:	dt	<=	138	;
						10'd518	:	dt	<=	157	;
						10'd519	:	dt	<=	177	;
						10'd520	:	dt	<=	175	;
						10'd521	:	dt	<=	171	;
						10'd522	:	dt	<=	152	;
						10'd523	:	dt	<=	114	;
						10'd524	:	dt	<=	112	;
						10'd525	:	dt	<=	163	;
						10'd526	:	dt	<=	175	;
						10'd527	:	dt	<=	177	;
						10'd528	:	dt	<=	178	;
						10'd529	:	dt	<=	180	;
						10'd530	:	dt	<=	180	;
						10'd531	:	dt	<=	181	;
						10'd532	:	dt	<=	106	;
						10'd533	:	dt	<=	108	;
						10'd534	:	dt	<=	94	;
						10'd535	:	dt	<=	95	;
						10'd536	:	dt	<=	79	;
						10'd537	:	dt	<=	38	;
						10'd538	:	dt	<=	62	;
						10'd539	:	dt	<=	87	;
						10'd540	:	dt	<=	131	;
						10'd541	:	dt	<=	159	;
						10'd542	:	dt	<=	140	;
						10'd543	:	dt	<=	124	;
						10'd544	:	dt	<=	128	;
						10'd545	:	dt	<=	142	;
						10'd546	:	dt	<=	162	;
						10'd547	:	dt	<=	181	;
						10'd548	:	dt	<=	180	;
						10'd549	:	dt	<=	166	;
						10'd550	:	dt	<=	146	;
						10'd551	:	dt	<=	112	;
						10'd552	:	dt	<=	110	;
						10'd553	:	dt	<=	162	;
						10'd554	:	dt	<=	175	;
						10'd555	:	dt	<=	177	;
						10'd556	:	dt	<=	179	;
						10'd557	:	dt	<=	180	;
						10'd558	:	dt	<=	181	;
						10'd559	:	dt	<=	182	;
						10'd560	:	dt	<=	107	;
						10'd561	:	dt	<=	108	;
						10'd562	:	dt	<=	93	;
						10'd563	:	dt	<=	97	;
						10'd564	:	dt	<=	74	;
						10'd565	:	dt	<=	38	;
						10'd566	:	dt	<=	64	;
						10'd567	:	dt	<=	86	;
						10'd568	:	dt	<=	118	;
						10'd569	:	dt	<=	155	;
						10'd570	:	dt	<=	147	;
						10'd571	:	dt	<=	129	;
						10'd572	:	dt	<=	127	;
						10'd573	:	dt	<=	145	;
						10'd574	:	dt	<=	164	;
						10'd575	:	dt	<=	182	;
						10'd576	:	dt	<=	181	;
						10'd577	:	dt	<=	162	;
						10'd578	:	dt	<=	137	;
						10'd579	:	dt	<=	104	;
						10'd580	:	dt	<=	111	;
						10'd581	:	dt	<=	164	;
						10'd582	:	dt	<=	175	;
						10'd583	:	dt	<=	177	;
						10'd584	:	dt	<=	179	;
						10'd585	:	dt	<=	181	;
						10'd586	:	dt	<=	182	;
						10'd587	:	dt	<=	182	;
						10'd588	:	dt	<=	108	;
						10'd589	:	dt	<=	109	;
						10'd590	:	dt	<=	93	;
						10'd591	:	dt	<=	100	;
						10'd592	:	dt	<=	70	;
						10'd593	:	dt	<=	39	;
						10'd594	:	dt	<=	66	;
						10'd595	:	dt	<=	86	;
						10'd596	:	dt	<=	108	;
						10'd597	:	dt	<=	147	;
						10'd598	:	dt	<=	154	;
						10'd599	:	dt	<=	137	;
						10'd600	:	dt	<=	128	;
						10'd601	:	dt	<=	141	;
						10'd602	:	dt	<=	161	;
						10'd603	:	dt	<=	179	;
						10'd604	:	dt	<=	177	;
						10'd605	:	dt	<=	157	;
						10'd606	:	dt	<=	132	;
						10'd607	:	dt	<=	100	;
						10'd608	:	dt	<=	113	;
						10'd609	:	dt	<=	165	;
						10'd610	:	dt	<=	175	;
						10'd611	:	dt	<=	177	;
						10'd612	:	dt	<=	179	;
						10'd613	:	dt	<=	181	;
						10'd614	:	dt	<=	182	;
						10'd615	:	dt	<=	182	;
						10'd616	:	dt	<=	111	;
						10'd617	:	dt	<=	111	;
						10'd618	:	dt	<=	93	;
						10'd619	:	dt	<=	103	;
						10'd620	:	dt	<=	66	;
						10'd621	:	dt	<=	40	;
						10'd622	:	dt	<=	68	;
						10'd623	:	dt	<=	86	;
						10'd624	:	dt	<=	102	;
						10'd625	:	dt	<=	136	;
						10'd626	:	dt	<=	156	;
						10'd627	:	dt	<=	145	;
						10'd628	:	dt	<=	134	;
						10'd629	:	dt	<=	136	;
						10'd630	:	dt	<=	155	;
						10'd631	:	dt	<=	174	;
						10'd632	:	dt	<=	169	;
						10'd633	:	dt	<=	150	;
						10'd634	:	dt	<=	128	;
						10'd635	:	dt	<=	98	;
						10'd636	:	dt	<=	113	;
						10'd637	:	dt	<=	166	;
						10'd638	:	dt	<=	176	;
						10'd639	:	dt	<=	178	;
						10'd640	:	dt	<=	180	;
						10'd641	:	dt	<=	181	;
						10'd642	:	dt	<=	182	;
						10'd643	:	dt	<=	182	;
						10'd644	:	dt	<=	114	;
						10'd645	:	dt	<=	113	;
						10'd646	:	dt	<=	95	;
						10'd647	:	dt	<=	107	;
						10'd648	:	dt	<=	62	;
						10'd649	:	dt	<=	41	;
						10'd650	:	dt	<=	69	;
						10'd651	:	dt	<=	85	;
						10'd652	:	dt	<=	98	;
						10'd653	:	dt	<=	121	;
						10'd654	:	dt	<=	149	;
						10'd655	:	dt	<=	151	;
						10'd656	:	dt	<=	143	;
						10'd657	:	dt	<=	137	;
						10'd658	:	dt	<=	149	;
						10'd659	:	dt	<=	166	;
						10'd660	:	dt	<=	161	;
						10'd661	:	dt	<=	143	;
						10'd662	:	dt	<=	122	;
						10'd663	:	dt	<=	95	;
						10'd664	:	dt	<=	117	;
						10'd665	:	dt	<=	167	;
						10'd666	:	dt	<=	176	;
						10'd667	:	dt	<=	178	;
						10'd668	:	dt	<=	180	;
						10'd669	:	dt	<=	181	;
						10'd670	:	dt	<=	181	;
						10'd671	:	dt	<=	182	;
						10'd672	:	dt	<=	118	;
						10'd673	:	dt	<=	114	;
						10'd674	:	dt	<=	97	;
						10'd675	:	dt	<=	108	;
						10'd676	:	dt	<=	57	;
						10'd677	:	dt	<=	42	;
						10'd678	:	dt	<=	68	;
						10'd679	:	dt	<=	84	;
						10'd680	:	dt	<=	95	;
						10'd681	:	dt	<=	110	;
						10'd682	:	dt	<=	135	;
						10'd683	:	dt	<=	151	;
						10'd684	:	dt	<=	149	;
						10'd685	:	dt	<=	142	;
						10'd686	:	dt	<=	141	;
						10'd687	:	dt	<=	151	;
						10'd688	:	dt	<=	152	;
						10'd689	:	dt	<=	136	;
						10'd690	:	dt	<=	117	;
						10'd691	:	dt	<=	95	;
						10'd692	:	dt	<=	126	;
						10'd693	:	dt	<=	168	;
						10'd694	:	dt	<=	174	;
						10'd695	:	dt	<=	176	;
						10'd696	:	dt	<=	178	;
						10'd697	:	dt	<=	178	;
						10'd698	:	dt	<=	180	;
						10'd699	:	dt	<=	180	;
						10'd700	:	dt	<=	120	;
						10'd701	:	dt	<=	113	;
						10'd702	:	dt	<=	98	;
						10'd703	:	dt	<=	108	;
						10'd704	:	dt	<=	52	;
						10'd705	:	dt	<=	43	;
						10'd706	:	dt	<=	67	;
						10'd707	:	dt	<=	82	;
						10'd708	:	dt	<=	93	;
						10'd709	:	dt	<=	105	;
						10'd710	:	dt	<=	121	;
						10'd711	:	dt	<=	147	;
						10'd712	:	dt	<=	151	;
						10'd713	:	dt	<=	143	;
						10'd714	:	dt	<=	133	;
						10'd715	:	dt	<=	135	;
						10'd716	:	dt	<=	139	;
						10'd717	:	dt	<=	126	;
						10'd718	:	dt	<=	111	;
						10'd719	:	dt	<=	99	;
						10'd720	:	dt	<=	139	;
						10'd721	:	dt	<=	169	;
						10'd722	:	dt	<=	173	;
						10'd723	:	dt	<=	174	;
						10'd724	:	dt	<=	176	;
						10'd725	:	dt	<=	177	;
						10'd726	:	dt	<=	178	;
						10'd727	:	dt	<=	179	;
						10'd728	:	dt	<=	122	;
						10'd729	:	dt	<=	112	;
						10'd730	:	dt	<=	100	;
						10'd731	:	dt	<=	107	;
						10'd732	:	dt	<=	47	;
						10'd733	:	dt	<=	43	;
						10'd734	:	dt	<=	66	;
						10'd735	:	dt	<=	79	;
						10'd736	:	dt	<=	90	;
						10'd737	:	dt	<=	102	;
						10'd738	:	dt	<=	113	;
						10'd739	:	dt	<=	140	;
						10'd740	:	dt	<=	149	;
						10'd741	:	dt	<=	138	;
						10'd742	:	dt	<=	128	;
						10'd743	:	dt	<=	127	;
						10'd744	:	dt	<=	126	;
						10'd745	:	dt	<=	119	;
						10'd746	:	dt	<=	107	;
						10'd747	:	dt	<=	100	;
						10'd748	:	dt	<=	146	;
						10'd749	:	dt	<=	168	;
						10'd750	:	dt	<=	170	;
						10'd751	:	dt	<=	173	;
						10'd752	:	dt	<=	175	;
						10'd753	:	dt	<=	176	;
						10'd754	:	dt	<=	178	;
						10'd755	:	dt	<=	178	;
						10'd756	:	dt	<=	123	;
						10'd757	:	dt	<=	110	;
						10'd758	:	dt	<=	101	;
						10'd759	:	dt	<=	105	;
						10'd760	:	dt	<=	45	;
						10'd761	:	dt	<=	45	;
						10'd762	:	dt	<=	64	;
						10'd763	:	dt	<=	74	;
						10'd764	:	dt	<=	85	;
						10'd765	:	dt	<=	97	;
						10'd766	:	dt	<=	108	;
						10'd767	:	dt	<=	134	;
						10'd768	:	dt	<=	145	;
						10'd769	:	dt	<=	133	;
						10'd770	:	dt	<=	128	;
						10'd771	:	dt	<=	129	;
						10'd772	:	dt	<=	125	;
						10'd773	:	dt	<=	117	;
						10'd774	:	dt	<=	103	;
						10'd775	:	dt	<=	98	;
						10'd776	:	dt	<=	147	;
						10'd777	:	dt	<=	166	;
						10'd778	:	dt	<=	168	;
						10'd779	:	dt	<=	171	;
						10'd780	:	dt	<=	173	;
						10'd781	:	dt	<=	175	;
						10'd782	:	dt	<=	176	;
						10'd783	:	dt	<=	176	;
					endcase
				end
				5'd2	:	begin
					case (cnt)
						10'd0	:	dt	<=	197	;
						10'd1	:	dt	<=	197	;
						10'd2	:	dt	<=	197	;
						10'd3	:	dt	<=	198	;
						10'd4	:	dt	<=	199	;
						10'd5	:	dt	<=	199	;
						10'd6	:	dt	<=	199	;
						10'd7	:	dt	<=	198	;
						10'd8	:	dt	<=	199	;
						10'd9	:	dt	<=	198	;
						10'd10	:	dt	<=	198	;
						10'd11	:	dt	<=	198	;
						10'd12	:	dt	<=	198	;
						10'd13	:	dt	<=	198	;
						10'd14	:	dt	<=	198	;
						10'd15	:	dt	<=	198	;
						10'd16	:	dt	<=	197	;
						10'd17	:	dt	<=	197	;
						10'd18	:	dt	<=	197	;
						10'd19	:	dt	<=	196	;
						10'd20	:	dt	<=	195	;
						10'd21	:	dt	<=	193	;
						10'd22	:	dt	<=	193	;
						10'd23	:	dt	<=	195	;
						10'd24	:	dt	<=	191	;
						10'd25	:	dt	<=	114	;
						10'd26	:	dt	<=	83	;
						10'd27	:	dt	<=	102	;
						10'd28	:	dt	<=	200	;
						10'd29	:	dt	<=	201	;
						10'd30	:	dt	<=	202	;
						10'd31	:	dt	<=	200	;
						10'd32	:	dt	<=	200	;
						10'd33	:	dt	<=	201	;
						10'd34	:	dt	<=	200	;
						10'd35	:	dt	<=	201	;
						10'd36	:	dt	<=	201	;
						10'd37	:	dt	<=	202	;
						10'd38	:	dt	<=	202	;
						10'd39	:	dt	<=	203	;
						10'd40	:	dt	<=	201	;
						10'd41	:	dt	<=	200	;
						10'd42	:	dt	<=	201	;
						10'd43	:	dt	<=	200	;
						10'd44	:	dt	<=	197	;
						10'd45	:	dt	<=	202	;
						10'd46	:	dt	<=	199	;
						10'd47	:	dt	<=	201	;
						10'd48	:	dt	<=	195	;
						10'd49	:	dt	<=	196	;
						10'd50	:	dt	<=	197	;
						10'd51	:	dt	<=	201	;
						10'd52	:	dt	<=	181	;
						10'd53	:	dt	<=	98	;
						10'd54	:	dt	<=	96	;
						10'd55	:	dt	<=	106	;
						10'd56	:	dt	<=	204	;
						10'd57	:	dt	<=	205	;
						10'd58	:	dt	<=	206	;
						10'd59	:	dt	<=	204	;
						10'd60	:	dt	<=	204	;
						10'd61	:	dt	<=	205	;
						10'd62	:	dt	<=	205	;
						10'd63	:	dt	<=	205	;
						10'd64	:	dt	<=	205	;
						10'd65	:	dt	<=	206	;
						10'd66	:	dt	<=	206	;
						10'd67	:	dt	<=	205	;
						10'd68	:	dt	<=	201	;
						10'd69	:	dt	<=	207	;
						10'd70	:	dt	<=	213	;
						10'd71	:	dt	<=	183	;
						10'd72	:	dt	<=	136	;
						10'd73	:	dt	<=	171	;
						10'd74	:	dt	<=	186	;
						10'd75	:	dt	<=	172	;
						10'd76	:	dt	<=	206	;
						10'd77	:	dt	<=	201	;
						10'd78	:	dt	<=	199	;
						10'd79	:	dt	<=	201	;
						10'd80	:	dt	<=	194	;
						10'd81	:	dt	<=	118	;
						10'd82	:	dt	<=	105	;
						10'd83	:	dt	<=	101	;
						10'd84	:	dt	<=	207	;
						10'd85	:	dt	<=	207	;
						10'd86	:	dt	<=	208	;
						10'd87	:	dt	<=	207	;
						10'd88	:	dt	<=	206	;
						10'd89	:	dt	<=	208	;
						10'd90	:	dt	<=	207	;
						10'd91	:	dt	<=	208	;
						10'd92	:	dt	<=	209	;
						10'd93	:	dt	<=	207	;
						10'd94	:	dt	<=	205	;
						10'd95	:	dt	<=	208	;
						10'd96	:	dt	<=	216	;
						10'd97	:	dt	<=	212	;
						10'd98	:	dt	<=	176	;
						10'd99	:	dt	<=	139	;
						10'd100	:	dt	<=	112	;
						10'd101	:	dt	<=	118	;
						10'd102	:	dt	<=	141	;
						10'd103	:	dt	<=	116	;
						10'd104	:	dt	<=	159	;
						10'd105	:	dt	<=	197	;
						10'd106	:	dt	<=	202	;
						10'd107	:	dt	<=	200	;
						10'd108	:	dt	<=	205	;
						10'd109	:	dt	<=	144	;
						10'd110	:	dt	<=	104	;
						10'd111	:	dt	<=	108	;
						10'd112	:	dt	<=	210	;
						10'd113	:	dt	<=	210	;
						10'd114	:	dt	<=	210	;
						10'd115	:	dt	<=	209	;
						10'd116	:	dt	<=	209	;
						10'd117	:	dt	<=	210	;
						10'd118	:	dt	<=	209	;
						10'd119	:	dt	<=	211	;
						10'd120	:	dt	<=	210	;
						10'd121	:	dt	<=	210	;
						10'd122	:	dt	<=	222	;
						10'd123	:	dt	<=	230	;
						10'd124	:	dt	<=	196	;
						10'd125	:	dt	<=	146	;
						10'd126	:	dt	<=	122	;
						10'd127	:	dt	<=	111	;
						10'd128	:	dt	<=	106	;
						10'd129	:	dt	<=	107	;
						10'd130	:	dt	<=	115	;
						10'd131	:	dt	<=	106	;
						10'd132	:	dt	<=	99	;
						10'd133	:	dt	<=	168	;
						10'd134	:	dt	<=	210	;
						10'd135	:	dt	<=	200	;
						10'd136	:	dt	<=	210	;
						10'd137	:	dt	<=	160	;
						10'd138	:	dt	<=	100	;
						10'd139	:	dt	<=	98	;
						10'd140	:	dt	<=	213	;
						10'd141	:	dt	<=	213	;
						10'd142	:	dt	<=	213	;
						10'd143	:	dt	<=	212	;
						10'd144	:	dt	<=	212	;
						10'd145	:	dt	<=	213	;
						10'd146	:	dt	<=	213	;
						10'd147	:	dt	<=	214	;
						10'd148	:	dt	<=	210	;
						10'd149	:	dt	<=	221	;
						10'd150	:	dt	<=	234	;
						10'd151	:	dt	<=	212	;
						10'd152	:	dt	<=	142	;
						10'd153	:	dt	<=	102	;
						10'd154	:	dt	<=	106	;
						10'd155	:	dt	<=	103	;
						10'd156	:	dt	<=	98	;
						10'd157	:	dt	<=	93	;
						10'd158	:	dt	<=	103	;
						10'd159	:	dt	<=	105	;
						10'd160	:	dt	<=	95	;
						10'd161	:	dt	<=	166	;
						10'd162	:	dt	<=	213	;
						10'd163	:	dt	<=	203	;
						10'd164	:	dt	<=	209	;
						10'd165	:	dt	<=	182	;
						10'd166	:	dt	<=	106	;
						10'd167	:	dt	<=	83	;
						10'd168	:	dt	<=	215	;
						10'd169	:	dt	<=	215	;
						10'd170	:	dt	<=	216	;
						10'd171	:	dt	<=	215	;
						10'd172	:	dt	<=	215	;
						10'd173	:	dt	<=	215	;
						10'd174	:	dt	<=	216	;
						10'd175	:	dt	<=	216	;
						10'd176	:	dt	<=	212	;
						10'd177	:	dt	<=	238	;
						10'd178	:	dt	<=	214	;
						10'd179	:	dt	<=	147	;
						10'd180	:	dt	<=	112	;
						10'd181	:	dt	<=	94	;
						10'd182	:	dt	<=	97	;
						10'd183	:	dt	<=	102	;
						10'd184	:	dt	<=	95	;
						10'd185	:	dt	<=	91	;
						10'd186	:	dt	<=	94	;
						10'd187	:	dt	<=	101	;
						10'd188	:	dt	<=	134	;
						10'd189	:	dt	<=	204	;
						10'd190	:	dt	<=	209	;
						10'd191	:	dt	<=	206	;
						10'd192	:	dt	<=	206	;
						10'd193	:	dt	<=	207	;
						10'd194	:	dt	<=	111	;
						10'd195	:	dt	<=	69	;
						10'd196	:	dt	<=	218	;
						10'd197	:	dt	<=	217	;
						10'd198	:	dt	<=	218	;
						10'd199	:	dt	<=	218	;
						10'd200	:	dt	<=	218	;
						10'd201	:	dt	<=	217	;
						10'd202	:	dt	<=	218	;
						10'd203	:	dt	<=	216	;
						10'd204	:	dt	<=	223	;
						10'd205	:	dt	<=	246	;
						10'd206	:	dt	<=	175	;
						10'd207	:	dt	<=	113	;
						10'd208	:	dt	<=	104	;
						10'd209	:	dt	<=	97	;
						10'd210	:	dt	<=	91	;
						10'd211	:	dt	<=	97	;
						10'd212	:	dt	<=	101	;
						10'd213	:	dt	<=	112	;
						10'd214	:	dt	<=	153	;
						10'd215	:	dt	<=	185	;
						10'd216	:	dt	<=	212	;
						10'd217	:	dt	<=	213	;
						10'd218	:	dt	<=	210	;
						10'd219	:	dt	<=	208	;
						10'd220	:	dt	<=	208	;
						10'd221	:	dt	<=	209	;
						10'd222	:	dt	<=	148	;
						10'd223	:	dt	<=	133	;
						10'd224	:	dt	<=	219	;
						10'd225	:	dt	<=	219	;
						10'd226	:	dt	<=	220	;
						10'd227	:	dt	<=	221	;
						10'd228	:	dt	<=	220	;
						10'd229	:	dt	<=	220	;
						10'd230	:	dt	<=	220	;
						10'd231	:	dt	<=	214	;
						10'd232	:	dt	<=	237	;
						10'd233	:	dt	<=	232	;
						10'd234	:	dt	<=	160	;
						10'd235	:	dt	<=	119	;
						10'd236	:	dt	<=	105	;
						10'd237	:	dt	<=	112	;
						10'd238	:	dt	<=	101	;
						10'd239	:	dt	<=	103	;
						10'd240	:	dt	<=	113	;
						10'd241	:	dt	<=	182	;
						10'd242	:	dt	<=	224	;
						10'd243	:	dt	<=	217	;
						10'd244	:	dt	<=	214	;
						10'd245	:	dt	<=	214	;
						10'd246	:	dt	<=	213	;
						10'd247	:	dt	<=	211	;
						10'd248	:	dt	<=	211	;
						10'd249	:	dt	<=	213	;
						10'd250	:	dt	<=	181	;
						10'd251	:	dt	<=	166	;
						10'd252	:	dt	<=	219	;
						10'd253	:	dt	<=	221	;
						10'd254	:	dt	<=	223	;
						10'd255	:	dt	<=	223	;
						10'd256	:	dt	<=	223	;
						10'd257	:	dt	<=	223	;
						10'd258	:	dt	<=	221	;
						10'd259	:	dt	<=	224	;
						10'd260	:	dt	<=	243	;
						10'd261	:	dt	<=	206	;
						10'd262	:	dt	<=	142	;
						10'd263	:	dt	<=	105	;
						10'd264	:	dt	<=	102	;
						10'd265	:	dt	<=	108	;
						10'd266	:	dt	<=	101	;
						10'd267	:	dt	<=	124	;
						10'd268	:	dt	<=	199	;
						10'd269	:	dt	<=	221	;
						10'd270	:	dt	<=	215	;
						10'd271	:	dt	<=	216	;
						10'd272	:	dt	<=	217	;
						10'd273	:	dt	<=	217	;
						10'd274	:	dt	<=	215	;
						10'd275	:	dt	<=	213	;
						10'd276	:	dt	<=	212	;
						10'd277	:	dt	<=	222	;
						10'd278	:	dt	<=	147	;
						10'd279	:	dt	<=	176	;
						10'd280	:	dt	<=	223	;
						10'd281	:	dt	<=	223	;
						10'd282	:	dt	<=	224	;
						10'd283	:	dt	<=	224	;
						10'd284	:	dt	<=	224	;
						10'd285	:	dt	<=	225	;
						10'd286	:	dt	<=	219	;
						10'd287	:	dt	<=	237	;
						10'd288	:	dt	<=	239	;
						10'd289	:	dt	<=	191	;
						10'd290	:	dt	<=	141	;
						10'd291	:	dt	<=	109	;
						10'd292	:	dt	<=	104	;
						10'd293	:	dt	<=	100	;
						10'd294	:	dt	<=	106	;
						10'd295	:	dt	<=	161	;
						10'd296	:	dt	<=	236	;
						10'd297	:	dt	<=	218	;
						10'd298	:	dt	<=	220	;
						10'd299	:	dt	<=	219	;
						10'd300	:	dt	<=	218	;
						10'd301	:	dt	<=	218	;
						10'd302	:	dt	<=	218	;
						10'd303	:	dt	<=	217	;
						10'd304	:	dt	<=	214	;
						10'd305	:	dt	<=	220	;
						10'd306	:	dt	<=	161	;
						10'd307	:	dt	<=	206	;
						10'd308	:	dt	<=	224	;
						10'd309	:	dt	<=	226	;
						10'd310	:	dt	<=	227	;
						10'd311	:	dt	<=	226	;
						10'd312	:	dt	<=	225	;
						10'd313	:	dt	<=	226	;
						10'd314	:	dt	<=	224	;
						10'd315	:	dt	<=	250	;
						10'd316	:	dt	<=	231	;
						10'd317	:	dt	<=	183	;
						10'd318	:	dt	<=	142	;
						10'd319	:	dt	<=	125	;
						10'd320	:	dt	<=	116	;
						10'd321	:	dt	<=	105	;
						10'd322	:	dt	<=	104	;
						10'd323	:	dt	<=	181	;
						10'd324	:	dt	<=	231	;
						10'd325	:	dt	<=	224	;
						10'd326	:	dt	<=	224	;
						10'd327	:	dt	<=	221	;
						10'd328	:	dt	<=	221	;
						10'd329	:	dt	<=	220	;
						10'd330	:	dt	<=	219	;
						10'd331	:	dt	<=	218	;
						10'd332	:	dt	<=	217	;
						10'd333	:	dt	<=	217	;
						10'd334	:	dt	<=	202	;
						10'd335	:	dt	<=	188	;
						10'd336	:	dt	<=	225	;
						10'd337	:	dt	<=	226	;
						10'd338	:	dt	<=	228	;
						10'd339	:	dt	<=	229	;
						10'd340	:	dt	<=	228	;
						10'd341	:	dt	<=	224	;
						10'd342	:	dt	<=	235	;
						10'd343	:	dt	<=	255	;
						10'd344	:	dt	<=	218	;
						10'd345	:	dt	<=	170	;
						10'd346	:	dt	<=	134	;
						10'd347	:	dt	<=	122	;
						10'd348	:	dt	<=	120	;
						10'd349	:	dt	<=	117	;
						10'd350	:	dt	<=	111	;
						10'd351	:	dt	<=	215	;
						10'd352	:	dt	<=	230	;
						10'd353	:	dt	<=	225	;
						10'd354	:	dt	<=	225	;
						10'd355	:	dt	<=	224	;
						10'd356	:	dt	<=	224	;
						10'd357	:	dt	<=	223	;
						10'd358	:	dt	<=	222	;
						10'd359	:	dt	<=	220	;
						10'd360	:	dt	<=	218	;
						10'd361	:	dt	<=	218	;
						10'd362	:	dt	<=	221	;
						10'd363	:	dt	<=	195	;
						10'd364	:	dt	<=	227	;
						10'd365	:	dt	<=	227	;
						10'd366	:	dt	<=	229	;
						10'd367	:	dt	<=	230	;
						10'd368	:	dt	<=	230	;
						10'd369	:	dt	<=	223	;
						10'd370	:	dt	<=	246	;
						10'd371	:	dt	<=	253	;
						10'd372	:	dt	<=	208	;
						10'd373	:	dt	<=	159	;
						10'd374	:	dt	<=	125	;
						10'd375	:	dt	<=	118	;
						10'd376	:	dt	<=	114	;
						10'd377	:	dt	<=	117	;
						10'd378	:	dt	<=	132	;
						10'd379	:	dt	<=	230	;
						10'd380	:	dt	<=	228	;
						10'd381	:	dt	<=	227	;
						10'd382	:	dt	<=	226	;
						10'd383	:	dt	<=	225	;
						10'd384	:	dt	<=	225	;
						10'd385	:	dt	<=	225	;
						10'd386	:	dt	<=	224	;
						10'd387	:	dt	<=	223	;
						10'd388	:	dt	<=	221	;
						10'd389	:	dt	<=	222	;
						10'd390	:	dt	<=	219	;
						10'd391	:	dt	<=	214	;
						10'd392	:	dt	<=	229	;
						10'd393	:	dt	<=	230	;
						10'd394	:	dt	<=	229	;
						10'd395	:	dt	<=	229	;
						10'd396	:	dt	<=	227	;
						10'd397	:	dt	<=	224	;
						10'd398	:	dt	<=	255	;
						10'd399	:	dt	<=	241	;
						10'd400	:	dt	<=	201	;
						10'd401	:	dt	<=	158	;
						10'd402	:	dt	<=	126	;
						10'd403	:	dt	<=	115	;
						10'd404	:	dt	<=	113	;
						10'd405	:	dt	<=	114	;
						10'd406	:	dt	<=	140	;
						10'd407	:	dt	<=	234	;
						10'd408	:	dt	<=	228	;
						10'd409	:	dt	<=	227	;
						10'd410	:	dt	<=	226	;
						10'd411	:	dt	<=	226	;
						10'd412	:	dt	<=	225	;
						10'd413	:	dt	<=	225	;
						10'd414	:	dt	<=	224	;
						10'd415	:	dt	<=	224	;
						10'd416	:	dt	<=	223	;
						10'd417	:	dt	<=	223	;
						10'd418	:	dt	<=	220	;
						10'd419	:	dt	<=	214	;
						10'd420	:	dt	<=	229	;
						10'd421	:	dt	<=	230	;
						10'd422	:	dt	<=	230	;
						10'd423	:	dt	<=	232	;
						10'd424	:	dt	<=	225	;
						10'd425	:	dt	<=	240	;
						10'd426	:	dt	<=	255	;
						10'd427	:	dt	<=	228	;
						10'd428	:	dt	<=	190	;
						10'd429	:	dt	<=	149	;
						10'd430	:	dt	<=	126	;
						10'd431	:	dt	<=	117	;
						10'd432	:	dt	<=	120	;
						10'd433	:	dt	<=	109	;
						10'd434	:	dt	<=	158	;
						10'd435	:	dt	<=	241	;
						10'd436	:	dt	<=	228	;
						10'd437	:	dt	<=	228	;
						10'd438	:	dt	<=	228	;
						10'd439	:	dt	<=	227	;
						10'd440	:	dt	<=	227	;
						10'd441	:	dt	<=	226	;
						10'd442	:	dt	<=	227	;
						10'd443	:	dt	<=	227	;
						10'd444	:	dt	<=	227	;
						10'd445	:	dt	<=	228	;
						10'd446	:	dt	<=	227	;
						10'd447	:	dt	<=	221	;
						10'd448	:	dt	<=	231	;
						10'd449	:	dt	<=	231	;
						10'd450	:	dt	<=	232	;
						10'd451	:	dt	<=	233	;
						10'd452	:	dt	<=	227	;
						10'd453	:	dt	<=	255	;
						10'd454	:	dt	<=	249	;
						10'd455	:	dt	<=	217	;
						10'd456	:	dt	<=	179	;
						10'd457	:	dt	<=	143	;
						10'd458	:	dt	<=	125	;
						10'd459	:	dt	<=	115	;
						10'd460	:	dt	<=	113	;
						10'd461	:	dt	<=	103	;
						10'd462	:	dt	<=	146	;
						10'd463	:	dt	<=	241	;
						10'd464	:	dt	<=	229	;
						10'd465	:	dt	<=	230	;
						10'd466	:	dt	<=	230	;
						10'd467	:	dt	<=	230	;
						10'd468	:	dt	<=	232	;
						10'd469	:	dt	<=	232	;
						10'd470	:	dt	<=	226	;
						10'd471	:	dt	<=	216	;
						10'd472	:	dt	<=	209	;
						10'd473	:	dt	<=	202	;
						10'd474	:	dt	<=	211	;
						10'd475	:	dt	<=	228	;
						10'd476	:	dt	<=	233	;
						10'd477	:	dt	<=	233	;
						10'd478	:	dt	<=	235	;
						10'd479	:	dt	<=	228	;
						10'd480	:	dt	<=	230	;
						10'd481	:	dt	<=	255	;
						10'd482	:	dt	<=	242	;
						10'd483	:	dt	<=	209	;
						10'd484	:	dt	<=	171	;
						10'd485	:	dt	<=	137	;
						10'd486	:	dt	<=	121	;
						10'd487	:	dt	<=	110	;
						10'd488	:	dt	<=	107	;
						10'd489	:	dt	<=	118	;
						10'd490	:	dt	<=	110	;
						10'd491	:	dt	<=	177	;
						10'd492	:	dt	<=	244	;
						10'd493	:	dt	<=	231	;
						10'd494	:	dt	<=	236	;
						10'd495	:	dt	<=	234	;
						10'd496	:	dt	<=	218	;
						10'd497	:	dt	<=	205	;
						10'd498	:	dt	<=	196	;
						10'd499	:	dt	<=	193	;
						10'd500	:	dt	<=	189	;
						10'd501	:	dt	<=	178	;
						10'd502	:	dt	<=	151	;
						10'd503	:	dt	<=	181	;
						10'd504	:	dt	<=	233	;
						10'd505	:	dt	<=	234	;
						10'd506	:	dt	<=	238	;
						10'd507	:	dt	<=	224	;
						10'd508	:	dt	<=	243	;
						10'd509	:	dt	<=	255	;
						10'd510	:	dt	<=	235	;
						10'd511	:	dt	<=	199	;
						10'd512	:	dt	<=	162	;
						10'd513	:	dt	<=	136	;
						10'd514	:	dt	<=	118	;
						10'd515	:	dt	<=	100	;
						10'd516	:	dt	<=	110	;
						10'd517	:	dt	<=	121	;
						10'd518	:	dt	<=	123	;
						10'd519	:	dt	<=	117	;
						10'd520	:	dt	<=	207	;
						10'd521	:	dt	<=	233	;
						10'd522	:	dt	<=	218	;
						10'd523	:	dt	<=	198	;
						10'd524	:	dt	<=	191	;
						10'd525	:	dt	<=	192	;
						10'd526	:	dt	<=	202	;
						10'd527	:	dt	<=	196	;
						10'd528	:	dt	<=	175	;
						10'd529	:	dt	<=	158	;
						10'd530	:	dt	<=	146	;
						10'd531	:	dt	<=	166	;
						10'd532	:	dt	<=	235	;
						10'd533	:	dt	<=	237	;
						10'd534	:	dt	<=	233	;
						10'd535	:	dt	<=	229	;
						10'd536	:	dt	<=	255	;
						10'd537	:	dt	<=	251	;
						10'd538	:	dt	<=	225	;
						10'd539	:	dt	<=	185	;
						10'd540	:	dt	<=	152	;
						10'd541	:	dt	<=	134	;
						10'd542	:	dt	<=	111	;
						10'd543	:	dt	<=	96	;
						10'd544	:	dt	<=	118	;
						10'd545	:	dt	<=	122	;
						10'd546	:	dt	<=	128	;
						10'd547	:	dt	<=	135	;
						10'd548	:	dt	<=	136	;
						10'd549	:	dt	<=	159	;
						10'd550	:	dt	<=	172	;
						10'd551	:	dt	<=	190	;
						10'd552	:	dt	<=	205	;
						10'd553	:	dt	<=	197	;
						10'd554	:	dt	<=	177	;
						10'd555	:	dt	<=	146	;
						10'd556	:	dt	<=	154	;
						10'd557	:	dt	<=	200	;
						10'd558	:	dt	<=	222	;
						10'd559	:	dt	<=	228	;
						10'd560	:	dt	<=	237	;
						10'd561	:	dt	<=	240	;
						10'd562	:	dt	<=	227	;
						10'd563	:	dt	<=	244	;
						10'd564	:	dt	<=	255	;
						10'd565	:	dt	<=	243	;
						10'd566	:	dt	<=	216	;
						10'd567	:	dt	<=	178	;
						10'd568	:	dt	<=	149	;
						10'd569	:	dt	<=	131	;
						10'd570	:	dt	<=	104	;
						10'd571	:	dt	<=	106	;
						10'd572	:	dt	<=	132	;
						10'd573	:	dt	<=	136	;
						10'd574	:	dt	<=	147	;
						10'd575	:	dt	<=	149	;
						10'd576	:	dt	<=	147	;
						10'd577	:	dt	<=	154	;
						10'd578	:	dt	<=	178	;
						10'd579	:	dt	<=	196	;
						10'd580	:	dt	<=	185	;
						10'd581	:	dt	<=	155	;
						10'd582	:	dt	<=	129	;
						10'd583	:	dt	<=	160	;
						10'd584	:	dt	<=	229	;
						10'd585	:	dt	<=	234	;
						10'd586	:	dt	<=	232	;
						10'd587	:	dt	<=	231	;
						10'd588	:	dt	<=	240	;
						10'd589	:	dt	<=	234	;
						10'd590	:	dt	<=	231	;
						10'd591	:	dt	<=	255	;
						10'd592	:	dt	<=	253	;
						10'd593	:	dt	<=	237	;
						10'd594	:	dt	<=	204	;
						10'd595	:	dt	<=	172	;
						10'd596	:	dt	<=	146	;
						10'd597	:	dt	<=	130	;
						10'd598	:	dt	<=	105	;
						10'd599	:	dt	<=	118	;
						10'd600	:	dt	<=	142	;
						10'd601	:	dt	<=	149	;
						10'd602	:	dt	<=	154	;
						10'd603	:	dt	<=	151	;
						10'd604	:	dt	<=	152	;
						10'd605	:	dt	<=	157	;
						10'd606	:	dt	<=	168	;
						10'd607	:	dt	<=	152	;
						10'd608	:	dt	<=	144	;
						10'd609	:	dt	<=	166	;
						10'd610	:	dt	<=	199	;
						10'd611	:	dt	<=	234	;
						10'd612	:	dt	<=	234	;
						10'd613	:	dt	<=	230	;
						10'd614	:	dt	<=	230	;
						10'd615	:	dt	<=	229	;
						10'd616	:	dt	<=	237	;
						10'd617	:	dt	<=	230	;
						10'd618	:	dt	<=	253	;
						10'd619	:	dt	<=	255	;
						10'd620	:	dt	<=	246	;
						10'd621	:	dt	<=	228	;
						10'd622	:	dt	<=	198	;
						10'd623	:	dt	<=	165	;
						10'd624	:	dt	<=	136	;
						10'd625	:	dt	<=	127	;
						10'd626	:	dt	<=	112	;
						10'd627	:	dt	<=	129	;
						10'd628	:	dt	<=	147	;
						10'd629	:	dt	<=	156	;
						10'd630	:	dt	<=	157	;
						10'd631	:	dt	<=	152	;
						10'd632	:	dt	<=	144	;
						10'd633	:	dt	<=	136	;
						10'd634	:	dt	<=	130	;
						10'd635	:	dt	<=	160	;
						10'd636	:	dt	<=	213	;
						10'd637	:	dt	<=	239	;
						10'd638	:	dt	<=	240	;
						10'd639	:	dt	<=	235	;
						10'd640	:	dt	<=	234	;
						10'd641	:	dt	<=	233	;
						10'd642	:	dt	<=	232	;
						10'd643	:	dt	<=	231	;
						10'd644	:	dt	<=	225	;
						10'd645	:	dt	<=	242	;
						10'd646	:	dt	<=	255	;
						10'd647	:	dt	<=	249	;
						10'd648	:	dt	<=	241	;
						10'd649	:	dt	<=	225	;
						10'd650	:	dt	<=	191	;
						10'd651	:	dt	<=	156	;
						10'd652	:	dt	<=	131	;
						10'd653	:	dt	<=	127	;
						10'd654	:	dt	<=	119	;
						10'd655	:	dt	<=	142	;
						10'd656	:	dt	<=	153	;
						10'd657	:	dt	<=	155	;
						10'd658	:	dt	<=	150	;
						10'd659	:	dt	<=	139	;
						10'd660	:	dt	<=	125	;
						10'd661	:	dt	<=	131	;
						10'd662	:	dt	<=	189	;
						10'd663	:	dt	<=	241	;
						10'd664	:	dt	<=	241	;
						10'd665	:	dt	<=	237	;
						10'd666	:	dt	<=	236	;
						10'd667	:	dt	<=	236	;
						10'd668	:	dt	<=	236	;
						10'd669	:	dt	<=	235	;
						10'd670	:	dt	<=	235	;
						10'd671	:	dt	<=	234	;
						10'd672	:	dt	<=	236	;
						10'd673	:	dt	<=	247	;
						10'd674	:	dt	<=	248	;
						10'd675	:	dt	<=	241	;
						10'd676	:	dt	<=	229	;
						10'd677	:	dt	<=	203	;
						10'd678	:	dt	<=	169	;
						10'd679	:	dt	<=	142	;
						10'd680	:	dt	<=	131	;
						10'd681	:	dt	<=	123	;
						10'd682	:	dt	<=	126	;
						10'd683	:	dt	<=	145	;
						10'd684	:	dt	<=	148	;
						10'd685	:	dt	<=	150	;
						10'd686	:	dt	<=	135	;
						10'd687	:	dt	<=	122	;
						10'd688	:	dt	<=	172	;
						10'd689	:	dt	<=	224	;
						10'd690	:	dt	<=	245	;
						10'd691	:	dt	<=	239	;
						10'd692	:	dt	<=	238	;
						10'd693	:	dt	<=	240	;
						10'd694	:	dt	<=	239	;
						10'd695	:	dt	<=	238	;
						10'd696	:	dt	<=	237	;
						10'd697	:	dt	<=	236	;
						10'd698	:	dt	<=	236	;
						10'd699	:	dt	<=	236	;
						10'd700	:	dt	<=	243	;
						10'd701	:	dt	<=	245	;
						10'd702	:	dt	<=	240	;
						10'd703	:	dt	<=	222	;
						10'd704	:	dt	<=	202	;
						10'd705	:	dt	<=	177	;
						10'd706	:	dt	<=	153	;
						10'd707	:	dt	<=	135	;
						10'd708	:	dt	<=	130	;
						10'd709	:	dt	<=	124	;
						10'd710	:	dt	<=	132	;
						10'd711	:	dt	<=	138	;
						10'd712	:	dt	<=	143	;
						10'd713	:	dt	<=	136	;
						10'd714	:	dt	<=	120	;
						10'd715	:	dt	<=	187	;
						10'd716	:	dt	<=	249	;
						10'd717	:	dt	<=	245	;
						10'd718	:	dt	<=	239	;
						10'd719	:	dt	<=	240	;
						10'd720	:	dt	<=	240	;
						10'd721	:	dt	<=	241	;
						10'd722	:	dt	<=	241	;
						10'd723	:	dt	<=	241	;
						10'd724	:	dt	<=	239	;
						10'd725	:	dt	<=	238	;
						10'd726	:	dt	<=	238	;
						10'd727	:	dt	<=	237	;
						10'd728	:	dt	<=	240	;
						10'd729	:	dt	<=	239	;
						10'd730	:	dt	<=	224	;
						10'd731	:	dt	<=	202	;
						10'd732	:	dt	<=	184	;
						10'd733	:	dt	<=	168	;
						10'd734	:	dt	<=	146	;
						10'd735	:	dt	<=	132	;
						10'd736	:	dt	<=	128	;
						10'd737	:	dt	<=	131	;
						10'd738	:	dt	<=	131	;
						10'd739	:	dt	<=	130	;
						10'd740	:	dt	<=	128	;
						10'd741	:	dt	<=	138	;
						10'd742	:	dt	<=	203	;
						10'd743	:	dt	<=	249	;
						10'd744	:	dt	<=	241	;
						10'd745	:	dt	<=	242	;
						10'd746	:	dt	<=	243	;
						10'd747	:	dt	<=	242	;
						10'd748	:	dt	<=	242	;
						10'd749	:	dt	<=	242	;
						10'd750	:	dt	<=	242	;
						10'd751	:	dt	<=	242	;
						10'd752	:	dt	<=	240	;
						10'd753	:	dt	<=	239	;
						10'd754	:	dt	<=	237	;
						10'd755	:	dt	<=	236	;
						10'd756	:	dt	<=	238	;
						10'd757	:	dt	<=	230	;
						10'd758	:	dt	<=	211	;
						10'd759	:	dt	<=	180	;
						10'd760	:	dt	<=	170	;
						10'd761	:	dt	<=	149	;
						10'd762	:	dt	<=	130	;
						10'd763	:	dt	<=	132	;
						10'd764	:	dt	<=	133	;
						10'd765	:	dt	<=	132	;
						10'd766	:	dt	<=	130	;
						10'd767	:	dt	<=	124	;
						10'd768	:	dt	<=	172	;
						10'd769	:	dt	<=	236	;
						10'd770	:	dt	<=	250	;
						10'd771	:	dt	<=	243	;
						10'd772	:	dt	<=	245	;
						10'd773	:	dt	<=	245	;
						10'd774	:	dt	<=	244	;
						10'd775	:	dt	<=	245	;
						10'd776	:	dt	<=	244	;
						10'd777	:	dt	<=	243	;
						10'd778	:	dt	<=	243	;
						10'd779	:	dt	<=	242	;
						10'd780	:	dt	<=	241	;
						10'd781	:	dt	<=	240	;
						10'd782	:	dt	<=	239	;
						10'd783	:	dt	<=	238	;
					endcase
				end
				5'd3	:	begin
					case (cnt)
						10'd0	:	dt	<=	188	;
						10'd1	:	dt	<=	191	;
						10'd2	:	dt	<=	193	;
						10'd3	:	dt	<=	195	;
						10'd4	:	dt	<=	199	;
						10'd5	:	dt	<=	201	;
						10'd6	:	dt	<=	202	;
						10'd7	:	dt	<=	203	;
						10'd8	:	dt	<=	203	;
						10'd9	:	dt	<=	203	;
						10'd10	:	dt	<=	204	;
						10'd11	:	dt	<=	204	;
						10'd12	:	dt	<=	204	;
						10'd13	:	dt	<=	203	;
						10'd14	:	dt	<=	202	;
						10'd15	:	dt	<=	198	;
						10'd16	:	dt	<=	216	;
						10'd17	:	dt	<=	217	;
						10'd18	:	dt	<=	135	;
						10'd19	:	dt	<=	181	;
						10'd20	:	dt	<=	200	;
						10'd21	:	dt	<=	195	;
						10'd22	:	dt	<=	194	;
						10'd23	:	dt	<=	193	;
						10'd24	:	dt	<=	190	;
						10'd25	:	dt	<=	189	;
						10'd26	:	dt	<=	187	;
						10'd27	:	dt	<=	185	;
						10'd28	:	dt	<=	190	;
						10'd29	:	dt	<=	194	;
						10'd30	:	dt	<=	196	;
						10'd31	:	dt	<=	197	;
						10'd32	:	dt	<=	200	;
						10'd33	:	dt	<=	202	;
						10'd34	:	dt	<=	204	;
						10'd35	:	dt	<=	206	;
						10'd36	:	dt	<=	207	;
						10'd37	:	dt	<=	207	;
						10'd38	:	dt	<=	206	;
						10'd39	:	dt	<=	205	;
						10'd40	:	dt	<=	206	;
						10'd41	:	dt	<=	206	;
						10'd42	:	dt	<=	205	;
						10'd43	:	dt	<=	200	;
						10'd44	:	dt	<=	220	;
						10'd45	:	dt	<=	206	;
						10'd46	:	dt	<=	122	;
						10'd47	:	dt	<=	155	;
						10'd48	:	dt	<=	207	;
						10'd49	:	dt	<=	196	;
						10'd50	:	dt	<=	195	;
						10'd51	:	dt	<=	195	;
						10'd52	:	dt	<=	193	;
						10'd53	:	dt	<=	191	;
						10'd54	:	dt	<=	188	;
						10'd55	:	dt	<=	187	;
						10'd56	:	dt	<=	192	;
						10'd57	:	dt	<=	195	;
						10'd58	:	dt	<=	198	;
						10'd59	:	dt	<=	199	;
						10'd60	:	dt	<=	203	;
						10'd61	:	dt	<=	205	;
						10'd62	:	dt	<=	206	;
						10'd63	:	dt	<=	208	;
						10'd64	:	dt	<=	209	;
						10'd65	:	dt	<=	209	;
						10'd66	:	dt	<=	209	;
						10'd67	:	dt	<=	208	;
						10'd68	:	dt	<=	208	;
						10'd69	:	dt	<=	207	;
						10'd70	:	dt	<=	207	;
						10'd71	:	dt	<=	202	;
						10'd72	:	dt	<=	219	;
						10'd73	:	dt	<=	195	;
						10'd74	:	dt	<=	123	;
						10'd75	:	dt	<=	146	;
						10'd76	:	dt	<=	209	;
						10'd77	:	dt	<=	197	;
						10'd78	:	dt	<=	197	;
						10'd79	:	dt	<=	197	;
						10'd80	:	dt	<=	195	;
						10'd81	:	dt	<=	191	;
						10'd82	:	dt	<=	190	;
						10'd83	:	dt	<=	188	;
						10'd84	:	dt	<=	193	;
						10'd85	:	dt	<=	197	;
						10'd86	:	dt	<=	200	;
						10'd87	:	dt	<=	201	;
						10'd88	:	dt	<=	204	;
						10'd89	:	dt	<=	207	;
						10'd90	:	dt	<=	209	;
						10'd91	:	dt	<=	210	;
						10'd92	:	dt	<=	211	;
						10'd93	:	dt	<=	211	;
						10'd94	:	dt	<=	211	;
						10'd95	:	dt	<=	210	;
						10'd96	:	dt	<=	210	;
						10'd97	:	dt	<=	209	;
						10'd98	:	dt	<=	208	;
						10'd99	:	dt	<=	205	;
						10'd100	:	dt	<=	219	;
						10'd101	:	dt	<=	197	;
						10'd102	:	dt	<=	123	;
						10'd103	:	dt	<=	142	;
						10'd104	:	dt	<=	209	;
						10'd105	:	dt	<=	199	;
						10'd106	:	dt	<=	200	;
						10'd107	:	dt	<=	197	;
						10'd108	:	dt	<=	195	;
						10'd109	:	dt	<=	194	;
						10'd110	:	dt	<=	192	;
						10'd111	:	dt	<=	190	;
						10'd112	:	dt	<=	196	;
						10'd113	:	dt	<=	199	;
						10'd114	:	dt	<=	202	;
						10'd115	:	dt	<=	204	;
						10'd116	:	dt	<=	206	;
						10'd117	:	dt	<=	209	;
						10'd118	:	dt	<=	211	;
						10'd119	:	dt	<=	212	;
						10'd120	:	dt	<=	213	;
						10'd121	:	dt	<=	213	;
						10'd122	:	dt	<=	213	;
						10'd123	:	dt	<=	212	;
						10'd124	:	dt	<=	212	;
						10'd125	:	dt	<=	212	;
						10'd126	:	dt	<=	210	;
						10'd127	:	dt	<=	206	;
						10'd128	:	dt	<=	223	;
						10'd129	:	dt	<=	221	;
						10'd130	:	dt	<=	143	;
						10'd131	:	dt	<=	135	;
						10'd132	:	dt	<=	207	;
						10'd133	:	dt	<=	202	;
						10'd134	:	dt	<=	201	;
						10'd135	:	dt	<=	200	;
						10'd136	:	dt	<=	197	;
						10'd137	:	dt	<=	196	;
						10'd138	:	dt	<=	194	;
						10'd139	:	dt	<=	191	;
						10'd140	:	dt	<=	199	;
						10'd141	:	dt	<=	201	;
						10'd142	:	dt	<=	203	;
						10'd143	:	dt	<=	207	;
						10'd144	:	dt	<=	209	;
						10'd145	:	dt	<=	211	;
						10'd146	:	dt	<=	213	;
						10'd147	:	dt	<=	215	;
						10'd148	:	dt	<=	216	;
						10'd149	:	dt	<=	216	;
						10'd150	:	dt	<=	216	;
						10'd151	:	dt	<=	216	;
						10'd152	:	dt	<=	215	;
						10'd153	:	dt	<=	213	;
						10'd154	:	dt	<=	212	;
						10'd155	:	dt	<=	207	;
						10'd156	:	dt	<=	229	;
						10'd157	:	dt	<=	225	;
						10'd158	:	dt	<=	143	;
						10'd159	:	dt	<=	127	;
						10'd160	:	dt	<=	206	;
						10'd161	:	dt	<=	203	;
						10'd162	:	dt	<=	202	;
						10'd163	:	dt	<=	201	;
						10'd164	:	dt	<=	198	;
						10'd165	:	dt	<=	196	;
						10'd166	:	dt	<=	195	;
						10'd167	:	dt	<=	193	;
						10'd168	:	dt	<=	199	;
						10'd169	:	dt	<=	203	;
						10'd170	:	dt	<=	206	;
						10'd171	:	dt	<=	209	;
						10'd172	:	dt	<=	212	;
						10'd173	:	dt	<=	214	;
						10'd174	:	dt	<=	216	;
						10'd175	:	dt	<=	217	;
						10'd176	:	dt	<=	218	;
						10'd177	:	dt	<=	218	;
						10'd178	:	dt	<=	218	;
						10'd179	:	dt	<=	217	;
						10'd180	:	dt	<=	216	;
						10'd181	:	dt	<=	216	;
						10'd182	:	dt	<=	215	;
						10'd183	:	dt	<=	208	;
						10'd184	:	dt	<=	234	;
						10'd185	:	dt	<=	215	;
						10'd186	:	dt	<=	133	;
						10'd187	:	dt	<=	125	;
						10'd188	:	dt	<=	209	;
						10'd189	:	dt	<=	205	;
						10'd190	:	dt	<=	203	;
						10'd191	:	dt	<=	202	;
						10'd192	:	dt	<=	200	;
						10'd193	:	dt	<=	197	;
						10'd194	:	dt	<=	196	;
						10'd195	:	dt	<=	195	;
						10'd196	:	dt	<=	201	;
						10'd197	:	dt	<=	205	;
						10'd198	:	dt	<=	209	;
						10'd199	:	dt	<=	211	;
						10'd200	:	dt	<=	215	;
						10'd201	:	dt	<=	217	;
						10'd202	:	dt	<=	219	;
						10'd203	:	dt	<=	220	;
						10'd204	:	dt	<=	221	;
						10'd205	:	dt	<=	220	;
						10'd206	:	dt	<=	220	;
						10'd207	:	dt	<=	220	;
						10'd208	:	dt	<=	218	;
						10'd209	:	dt	<=	218	;
						10'd210	:	dt	<=	217	;
						10'd211	:	dt	<=	210	;
						10'd212	:	dt	<=	234	;
						10'd213	:	dt	<=	214	;
						10'd214	:	dt	<=	136	;
						10'd215	:	dt	<=	127	;
						10'd216	:	dt	<=	212	;
						10'd217	:	dt	<=	208	;
						10'd218	:	dt	<=	206	;
						10'd219	:	dt	<=	204	;
						10'd220	:	dt	<=	202	;
						10'd221	:	dt	<=	199	;
						10'd222	:	dt	<=	197	;
						10'd223	:	dt	<=	196	;
						10'd224	:	dt	<=	203	;
						10'd225	:	dt	<=	207	;
						10'd226	:	dt	<=	211	;
						10'd227	:	dt	<=	215	;
						10'd228	:	dt	<=	217	;
						10'd229	:	dt	<=	218	;
						10'd230	:	dt	<=	221	;
						10'd231	:	dt	<=	222	;
						10'd232	:	dt	<=	223	;
						10'd233	:	dt	<=	223	;
						10'd234	:	dt	<=	223	;
						10'd235	:	dt	<=	223	;
						10'd236	:	dt	<=	222	;
						10'd237	:	dt	<=	220	;
						10'd238	:	dt	<=	219	;
						10'd239	:	dt	<=	215	;
						10'd240	:	dt	<=	245	;
						10'd241	:	dt	<=	211	;
						10'd242	:	dt	<=	138	;
						10'd243	:	dt	<=	127	;
						10'd244	:	dt	<=	212	;
						10'd245	:	dt	<=	209	;
						10'd246	:	dt	<=	208	;
						10'd247	:	dt	<=	206	;
						10'd248	:	dt	<=	204	;
						10'd249	:	dt	<=	201	;
						10'd250	:	dt	<=	200	;
						10'd251	:	dt	<=	197	;
						10'd252	:	dt	<=	205	;
						10'd253	:	dt	<=	209	;
						10'd254	:	dt	<=	213	;
						10'd255	:	dt	<=	216	;
						10'd256	:	dt	<=	218	;
						10'd257	:	dt	<=	221	;
						10'd258	:	dt	<=	223	;
						10'd259	:	dt	<=	225	;
						10'd260	:	dt	<=	225	;
						10'd261	:	dt	<=	226	;
						10'd262	:	dt	<=	225	;
						10'd263	:	dt	<=	225	;
						10'd264	:	dt	<=	224	;
						10'd265	:	dt	<=	221	;
						10'd266	:	dt	<=	222	;
						10'd267	:	dt	<=	211	;
						10'd268	:	dt	<=	196	;
						10'd269	:	dt	<=	171	;
						10'd270	:	dt	<=	117	;
						10'd271	:	dt	<=	125	;
						10'd272	:	dt	<=	218	;
						10'd273	:	dt	<=	209	;
						10'd274	:	dt	<=	209	;
						10'd275	:	dt	<=	208	;
						10'd276	:	dt	<=	205	;
						10'd277	:	dt	<=	202	;
						10'd278	:	dt	<=	199	;
						10'd279	:	dt	<=	197	;
						10'd280	:	dt	<=	206	;
						10'd281	:	dt	<=	211	;
						10'd282	:	dt	<=	215	;
						10'd283	:	dt	<=	218	;
						10'd284	:	dt	<=	221	;
						10'd285	:	dt	<=	224	;
						10'd286	:	dt	<=	226	;
						10'd287	:	dt	<=	227	;
						10'd288	:	dt	<=	228	;
						10'd289	:	dt	<=	228	;
						10'd290	:	dt	<=	228	;
						10'd291	:	dt	<=	227	;
						10'd292	:	dt	<=	225	;
						10'd293	:	dt	<=	228	;
						10'd294	:	dt	<=	248	;
						10'd295	:	dt	<=	205	;
						10'd296	:	dt	<=	135	;
						10'd297	:	dt	<=	103	;
						10'd298	:	dt	<=	83	;
						10'd299	:	dt	<=	146	;
						10'd300	:	dt	<=	224	;
						10'd301	:	dt	<=	210	;
						10'd302	:	dt	<=	211	;
						10'd303	:	dt	<=	210	;
						10'd304	:	dt	<=	206	;
						10'd305	:	dt	<=	204	;
						10'd306	:	dt	<=	201	;
						10'd307	:	dt	<=	199	;
						10'd308	:	dt	<=	208	;
						10'd309	:	dt	<=	213	;
						10'd310	:	dt	<=	217	;
						10'd311	:	dt	<=	220	;
						10'd312	:	dt	<=	224	;
						10'd313	:	dt	<=	226	;
						10'd314	:	dt	<=	227	;
						10'd315	:	dt	<=	229	;
						10'd316	:	dt	<=	230	;
						10'd317	:	dt	<=	230	;
						10'd318	:	dt	<=	229	;
						10'd319	:	dt	<=	226	;
						10'd320	:	dt	<=	224	;
						10'd321	:	dt	<=	206	;
						10'd322	:	dt	<=	203	;
						10'd323	:	dt	<=	208	;
						10'd324	:	dt	<=	162	;
						10'd325	:	dt	<=	122	;
						10'd326	:	dt	<=	67	;
						10'd327	:	dt	<=	188	;
						10'd328	:	dt	<=	226	;
						10'd329	:	dt	<=	212	;
						10'd330	:	dt	<=	214	;
						10'd331	:	dt	<=	212	;
						10'd332	:	dt	<=	209	;
						10'd333	:	dt	<=	206	;
						10'd334	:	dt	<=	203	;
						10'd335	:	dt	<=	201	;
						10'd336	:	dt	<=	210	;
						10'd337	:	dt	<=	214	;
						10'd338	:	dt	<=	218	;
						10'd339	:	dt	<=	222	;
						10'd340	:	dt	<=	225	;
						10'd341	:	dt	<=	227	;
						10'd342	:	dt	<=	230	;
						10'd343	:	dt	<=	230	;
						10'd344	:	dt	<=	232	;
						10'd345	:	dt	<=	232	;
						10'd346	:	dt	<=	226	;
						10'd347	:	dt	<=	241	;
						10'd348	:	dt	<=	241	;
						10'd349	:	dt	<=	173	;
						10'd350	:	dt	<=	112	;
						10'd351	:	dt	<=	174	;
						10'd352	:	dt	<=	233	;
						10'd353	:	dt	<=	151	;
						10'd354	:	dt	<=	109	;
						10'd355	:	dt	<=	168	;
						10'd356	:	dt	<=	210	;
						10'd357	:	dt	<=	221	;
						10'd358	:	dt	<=	216	;
						10'd359	:	dt	<=	213	;
						10'd360	:	dt	<=	210	;
						10'd361	:	dt	<=	208	;
						10'd362	:	dt	<=	205	;
						10'd363	:	dt	<=	203	;
						10'd364	:	dt	<=	210	;
						10'd365	:	dt	<=	216	;
						10'd366	:	dt	<=	219	;
						10'd367	:	dt	<=	223	;
						10'd368	:	dt	<=	226	;
						10'd369	:	dt	<=	229	;
						10'd370	:	dt	<=	231	;
						10'd371	:	dt	<=	233	;
						10'd372	:	dt	<=	228	;
						10'd373	:	dt	<=	236	;
						10'd374	:	dt	<=	199	;
						10'd375	:	dt	<=	159	;
						10'd376	:	dt	<=	215	;
						10'd377	:	dt	<=	180	;
						10'd378	:	dt	<=	130	;
						10'd379	:	dt	<=	150	;
						10'd380	:	dt	<=	240	;
						10'd381	:	dt	<=	144	;
						10'd382	:	dt	<=	123	;
						10'd383	:	dt	<=	104	;
						10'd384	:	dt	<=	137	;
						10'd385	:	dt	<=	161	;
						10'd386	:	dt	<=	215	;
						10'd387	:	dt	<=	215	;
						10'd388	:	dt	<=	211	;
						10'd389	:	dt	<=	210	;
						10'd390	:	dt	<=	208	;
						10'd391	:	dt	<=	205	;
						10'd392	:	dt	<=	211	;
						10'd393	:	dt	<=	217	;
						10'd394	:	dt	<=	221	;
						10'd395	:	dt	<=	224	;
						10'd396	:	dt	<=	228	;
						10'd397	:	dt	<=	231	;
						10'd398	:	dt	<=	232	;
						10'd399	:	dt	<=	232	;
						10'd400	:	dt	<=	247	;
						10'd401	:	dt	<=	248	;
						10'd402	:	dt	<=	200	;
						10'd403	:	dt	<=	135	;
						10'd404	:	dt	<=	166	;
						10'd405	:	dt	<=	204	;
						10'd406	:	dt	<=	149	;
						10'd407	:	dt	<=	127	;
						10'd408	:	dt	<=	202	;
						10'd409	:	dt	<=	154	;
						10'd410	:	dt	<=	142	;
						10'd411	:	dt	<=	123	;
						10'd412	:	dt	<=	154	;
						10'd413	:	dt	<=	116	;
						10'd414	:	dt	<=	187	;
						10'd415	:	dt	<=	223	;
						10'd416	:	dt	<=	211	;
						10'd417	:	dt	<=	211	;
						10'd418	:	dt	<=	209	;
						10'd419	:	dt	<=	207	;
						10'd420	:	dt	<=	213	;
						10'd421	:	dt	<=	218	;
						10'd422	:	dt	<=	222	;
						10'd423	:	dt	<=	226	;
						10'd424	:	dt	<=	229	;
						10'd425	:	dt	<=	232	;
						10'd426	:	dt	<=	232	;
						10'd427	:	dt	<=	240	;
						10'd428	:	dt	<=	251	;
						10'd429	:	dt	<=	234	;
						10'd430	:	dt	<=	220	;
						10'd431	:	dt	<=	177	;
						10'd432	:	dt	<=	135	;
						10'd433	:	dt	<=	198	;
						10'd434	:	dt	<=	148	;
						10'd435	:	dt	<=	114	;
						10'd436	:	dt	<=	166	;
						10'd437	:	dt	<=	166	;
						10'd438	:	dt	<=	154	;
						10'd439	:	dt	<=	134	;
						10'd440	:	dt	<=	149	;
						10'd441	:	dt	<=	103	;
						10'd442	:	dt	<=	177	;
						10'd443	:	dt	<=	226	;
						10'd444	:	dt	<=	213	;
						10'd445	:	dt	<=	213	;
						10'd446	:	dt	<=	210	;
						10'd447	:	dt	<=	208	;
						10'd448	:	dt	<=	212	;
						10'd449	:	dt	<=	218	;
						10'd450	:	dt	<=	223	;
						10'd451	:	dt	<=	226	;
						10'd452	:	dt	<=	230	;
						10'd453	:	dt	<=	233	;
						10'd454	:	dt	<=	232	;
						10'd455	:	dt	<=	255	;
						10'd456	:	dt	<=	250	;
						10'd457	:	dt	<=	221	;
						10'd458	:	dt	<=	229	;
						10'd459	:	dt	<=	182	;
						10'd460	:	dt	<=	128	;
						10'd461	:	dt	<=	167	;
						10'd462	:	dt	<=	147	;
						10'd463	:	dt	<=	113	;
						10'd464	:	dt	<=	156	;
						10'd465	:	dt	<=	127	;
						10'd466	:	dt	<=	118	;
						10'd467	:	dt	<=	148	;
						10'd468	:	dt	<=	127	;
						10'd469	:	dt	<=	93	;
						10'd470	:	dt	<=	174	;
						10'd471	:	dt	<=	229	;
						10'd472	:	dt	<=	214	;
						10'd473	:	dt	<=	215	;
						10'd474	:	dt	<=	212	;
						10'd475	:	dt	<=	210	;
						10'd476	:	dt	<=	212	;
						10'd477	:	dt	<=	217	;
						10'd478	:	dt	<=	223	;
						10'd479	:	dt	<=	226	;
						10'd480	:	dt	<=	230	;
						10'd481	:	dt	<=	232	;
						10'd482	:	dt	<=	232	;
						10'd483	:	dt	<=	249	;
						10'd484	:	dt	<=	242	;
						10'd485	:	dt	<=	194	;
						10'd486	:	dt	<=	200	;
						10'd487	:	dt	<=	180	;
						10'd488	:	dt	<=	120	;
						10'd489	:	dt	<=	134	;
						10'd490	:	dt	<=	144	;
						10'd491	:	dt	<=	96	;
						10'd492	:	dt	<=	185	;
						10'd493	:	dt	<=	187	;
						10'd494	:	dt	<=	100	;
						10'd495	:	dt	<=	170	;
						10'd496	:	dt	<=	156	;
						10'd497	:	dt	<=	95	;
						10'd498	:	dt	<=	150	;
						10'd499	:	dt	<=	230	;
						10'd500	:	dt	<=	214	;
						10'd501	:	dt	<=	213	;
						10'd502	:	dt	<=	211	;
						10'd503	:	dt	<=	209	;
						10'd504	:	dt	<=	215	;
						10'd505	:	dt	<=	219	;
						10'd506	:	dt	<=	224	;
						10'd507	:	dt	<=	229	;
						10'd508	:	dt	<=	231	;
						10'd509	:	dt	<=	234	;
						10'd510	:	dt	<=	236	;
						10'd511	:	dt	<=	238	;
						10'd512	:	dt	<=	238	;
						10'd513	:	dt	<=	212	;
						10'd514	:	dt	<=	199	;
						10'd515	:	dt	<=	159	;
						10'd516	:	dt	<=	99	;
						10'd517	:	dt	<=	128	;
						10'd518	:	dt	<=	128	;
						10'd519	:	dt	<=	77	;
						10'd520	:	dt	<=	180	;
						10'd521	:	dt	<=	194	;
						10'd522	:	dt	<=	104	;
						10'd523	:	dt	<=	152	;
						10'd524	:	dt	<=	162	;
						10'd525	:	dt	<=	92	;
						10'd526	:	dt	<=	130	;
						10'd527	:	dt	<=	230	;
						10'd528	:	dt	<=	215	;
						10'd529	:	dt	<=	214	;
						10'd530	:	dt	<=	210	;
						10'd531	:	dt	<=	207	;
						10'd532	:	dt	<=	215	;
						10'd533	:	dt	<=	220	;
						10'd534	:	dt	<=	225	;
						10'd535	:	dt	<=	228	;
						10'd536	:	dt	<=	231	;
						10'd537	:	dt	<=	234	;
						10'd538	:	dt	<=	236	;
						10'd539	:	dt	<=	242	;
						10'd540	:	dt	<=	251	;
						10'd541	:	dt	<=	233	;
						10'd542	:	dt	<=	211	;
						10'd543	:	dt	<=	148	;
						10'd544	:	dt	<=	123	;
						10'd545	:	dt	<=	132	;
						10'd546	:	dt	<=	141	;
						10'd547	:	dt	<=	105	;
						10'd548	:	dt	<=	164	;
						10'd549	:	dt	<=	168	;
						10'd550	:	dt	<=	143	;
						10'd551	:	dt	<=	145	;
						10'd552	:	dt	<=	133	;
						10'd553	:	dt	<=	87	;
						10'd554	:	dt	<=	174	;
						10'd555	:	dt	<=	227	;
						10'd556	:	dt	<=	213	;
						10'd557	:	dt	<=	214	;
						10'd558	:	dt	<=	215	;
						10'd559	:	dt	<=	218	;
						10'd560	:	dt	<=	214	;
						10'd561	:	dt	<=	220	;
						10'd562	:	dt	<=	226	;
						10'd563	:	dt	<=	229	;
						10'd564	:	dt	<=	231	;
						10'd565	:	dt	<=	234	;
						10'd566	:	dt	<=	235	;
						10'd567	:	dt	<=	240	;
						10'd568	:	dt	<=	255	;
						10'd569	:	dt	<=	240	;
						10'd570	:	dt	<=	226	;
						10'd571	:	dt	<=	153	;
						10'd572	:	dt	<=	131	;
						10'd573	:	dt	<=	131	;
						10'd574	:	dt	<=	155	;
						10'd575	:	dt	<=	168	;
						10'd576	:	dt	<=	220	;
						10'd577	:	dt	<=	197	;
						10'd578	:	dt	<=	168	;
						10'd579	:	dt	<=	147	;
						10'd580	:	dt	<=	97	;
						10'd581	:	dt	<=	115	;
						10'd582	:	dt	<=	229	;
						10'd583	:	dt	<=	227	;
						10'd584	:	dt	<=	228	;
						10'd585	:	dt	<=	225	;
						10'd586	:	dt	<=	204	;
						10'd587	:	dt	<=	161	;
						10'd588	:	dt	<=	217	;
						10'd589	:	dt	<=	223	;
						10'd590	:	dt	<=	229	;
						10'd591	:	dt	<=	233	;
						10'd592	:	dt	<=	235	;
						10'd593	:	dt	<=	238	;
						10'd594	:	dt	<=	241	;
						10'd595	:	dt	<=	243	;
						10'd596	:	dt	<=	255	;
						10'd597	:	dt	<=	249	;
						10'd598	:	dt	<=	221	;
						10'd599	:	dt	<=	169	;
						10'd600	:	dt	<=	150	;
						10'd601	:	dt	<=	139	;
						10'd602	:	dt	<=	203	;
						10'd603	:	dt	<=	232	;
						10'd604	:	dt	<=	209	;
						10'd605	:	dt	<=	176	;
						10'd606	:	dt	<=	139	;
						10'd607	:	dt	<=	131	;
						10'd608	:	dt	<=	93	;
						10'd609	:	dt	<=	182	;
						10'd610	:	dt	<=	234	;
						10'd611	:	dt	<=	193	;
						10'd612	:	dt	<=	166	;
						10'd613	:	dt	<=	138	;
						10'd614	:	dt	<=	92	;
						10'd615	:	dt	<=	66	;
						10'd616	:	dt	<=	165	;
						10'd617	:	dt	<=	165	;
						10'd618	:	dt	<=	167	;
						10'd619	:	dt	<=	169	;
						10'd620	:	dt	<=	170	;
						10'd621	:	dt	<=	170	;
						10'd622	:	dt	<=	167	;
						10'd623	:	dt	<=	167	;
						10'd624	:	dt	<=	238	;
						10'd625	:	dt	<=	245	;
						10'd626	:	dt	<=	212	;
						10'd627	:	dt	<=	191	;
						10'd628	:	dt	<=	163	;
						10'd629	:	dt	<=	154	;
						10'd630	:	dt	<=	214	;
						10'd631	:	dt	<=	223	;
						10'd632	:	dt	<=	188	;
						10'd633	:	dt	<=	155	;
						10'd634	:	dt	<=	131	;
						10'd635	:	dt	<=	118	;
						10'd636	:	dt	<=	95	;
						10'd637	:	dt	<=	124	;
						10'd638	:	dt	<=	103	;
						10'd639	:	dt	<=	65	;
						10'd640	:	dt	<=	50	;
						10'd641	:	dt	<=	47	;
						10'd642	:	dt	<=	54	;
						10'd643	:	dt	<=	59	;
						10'd644	:	dt	<=	139	;
						10'd645	:	dt	<=	141	;
						10'd646	:	dt	<=	140	;
						10'd647	:	dt	<=	141	;
						10'd648	:	dt	<=	140	;
						10'd649	:	dt	<=	137	;
						10'd650	:	dt	<=	140	;
						10'd651	:	dt	<=	124	;
						10'd652	:	dt	<=	201	;
						10'd653	:	dt	<=	244	;
						10'd654	:	dt	<=	213	;
						10'd655	:	dt	<=	195	;
						10'd656	:	dt	<=	177	;
						10'd657	:	dt	<=	145	;
						10'd658	:	dt	<=	180	;
						10'd659	:	dt	<=	191	;
						10'd660	:	dt	<=	162	;
						10'd661	:	dt	<=	136	;
						10'd662	:	dt	<=	120	;
						10'd663	:	dt	<=	100	;
						10'd664	:	dt	<=	70	;
						10'd665	:	dt	<=	49	;
						10'd666	:	dt	<=	47	;
						10'd667	:	dt	<=	50	;
						10'd668	:	dt	<=	57	;
						10'd669	:	dt	<=	54	;
						10'd670	:	dt	<=	47	;
						10'd671	:	dt	<=	50	;
						10'd672	:	dt	<=	147	;
						10'd673	:	dt	<=	148	;
						10'd674	:	dt	<=	147	;
						10'd675	:	dt	<=	147	;
						10'd676	:	dt	<=	147	;
						10'd677	:	dt	<=	148	;
						10'd678	:	dt	<=	158	;
						10'd679	:	dt	<=	126	;
						10'd680	:	dt	<=	124	;
						10'd681	:	dt	<=	242	;
						10'd682	:	dt	<=	215	;
						10'd683	:	dt	<=	194	;
						10'd684	:	dt	<=	176	;
						10'd685	:	dt	<=	136	;
						10'd686	:	dt	<=	137	;
						10'd687	:	dt	<=	135	;
						10'd688	:	dt	<=	129	;
						10'd689	:	dt	<=	115	;
						10'd690	:	dt	<=	100	;
						10'd691	:	dt	<=	70	;
						10'd692	:	dt	<=	53	;
						10'd693	:	dt	<=	56	;
						10'd694	:	dt	<=	57	;
						10'd695	:	dt	<=	49	;
						10'd696	:	dt	<=	48	;
						10'd697	:	dt	<=	58	;
						10'd698	:	dt	<=	53	;
						10'd699	:	dt	<=	46	;
						10'd700	:	dt	<=	148	;
						10'd701	:	dt	<=	148	;
						10'd702	:	dt	<=	146	;
						10'd703	:	dt	<=	146	;
						10'd704	:	dt	<=	146	;
						10'd705	:	dt	<=	146	;
						10'd706	:	dt	<=	148	;
						10'd707	:	dt	<=	121	;
						10'd708	:	dt	<=	64	;
						10'd709	:	dt	<=	148	;
						10'd710	:	dt	<=	207	;
						10'd711	:	dt	<=	197	;
						10'd712	:	dt	<=	154	;
						10'd713	:	dt	<=	117	;
						10'd714	:	dt	<=	119	;
						10'd715	:	dt	<=	116	;
						10'd716	:	dt	<=	119	;
						10'd717	:	dt	<=	91	;
						10'd718	:	dt	<=	54	;
						10'd719	:	dt	<=	69	;
						10'd720	:	dt	<=	46	;
						10'd721	:	dt	<=	43	;
						10'd722	:	dt	<=	53	;
						10'd723	:	dt	<=	52	;
						10'd724	:	dt	<=	44	;
						10'd725	:	dt	<=	48	;
						10'd726	:	dt	<=	56	;
						10'd727	:	dt	<=	55	;
						10'd728	:	dt	<=	148	;
						10'd729	:	dt	<=	150	;
						10'd730	:	dt	<=	151	;
						10'd731	:	dt	<=	149	;
						10'd732	:	dt	<=	148	;
						10'd733	:	dt	<=	149	;
						10'd734	:	dt	<=	143	;
						10'd735	:	dt	<=	95	;
						10'd736	:	dt	<=	79	;
						10'd737	:	dt	<=	74	;
						10'd738	:	dt	<=	115	;
						10'd739	:	dt	<=	144	;
						10'd740	:	dt	<=	125	;
						10'd741	:	dt	<=	120	;
						10'd742	:	dt	<=	112	;
						10'd743	:	dt	<=	105	;
						10'd744	:	dt	<=	93	;
						10'd745	:	dt	<=	52	;
						10'd746	:	dt	<=	24	;
						10'd747	:	dt	<=	53	;
						10'd748	:	dt	<=	63	;
						10'd749	:	dt	<=	33	;
						10'd750	:	dt	<=	41	;
						10'd751	:	dt	<=	51	;
						10'd752	:	dt	<=	48	;
						10'd753	:	dt	<=	45	;
						10'd754	:	dt	<=	49	;
						10'd755	:	dt	<=	55	;
						10'd756	:	dt	<=	149	;
						10'd757	:	dt	<=	150	;
						10'd758	:	dt	<=	150	;
						10'd759	:	dt	<=	148	;
						10'd760	:	dt	<=	147	;
						10'd761	:	dt	<=	151	;
						10'd762	:	dt	<=	124	;
						10'd763	:	dt	<=	82	;
						10'd764	:	dt	<=	84	;
						10'd765	:	dt	<=	81	;
						10'd766	:	dt	<=	69	;
						10'd767	:	dt	<=	81	;
						10'd768	:	dt	<=	111	;
						10'd769	:	dt	<=	103	;
						10'd770	:	dt	<=	84	;
						10'd771	:	dt	<=	75	;
						10'd772	:	dt	<=	53	;
						10'd773	:	dt	<=	28	;
						10'd774	:	dt	<=	26	;
						10'd775	:	dt	<=	40	;
						10'd776	:	dt	<=	64	;
						10'd777	:	dt	<=	48	;
						10'd778	:	dt	<=	29	;
						10'd779	:	dt	<=	46	;
						10'd780	:	dt	<=	49	;
						10'd781	:	dt	<=	46	;
						10'd782	:	dt	<=	46	;
						10'd783	:	dt	<=	53	;
					endcase
				end
				5'd4	:	begin
					case (cnt)
						10'd0	:	dt	<=	191	;
						10'd1	:	dt	<=	192	;
						10'd2	:	dt	<=	192	;
						10'd3	:	dt	<=	192	;
						10'd4	:	dt	<=	192	;
						10'd5	:	dt	<=	193	;
						10'd6	:	dt	<=	193	;
						10'd7	:	dt	<=	193	;
						10'd8	:	dt	<=	193	;
						10'd9	:	dt	<=	192	;
						10'd10	:	dt	<=	193	;
						10'd11	:	dt	<=	193	;
						10'd12	:	dt	<=	192	;
						10'd13	:	dt	<=	192	;
						10'd14	:	dt	<=	192	;
						10'd15	:	dt	<=	191	;
						10'd16	:	dt	<=	190	;
						10'd17	:	dt	<=	187	;
						10'd18	:	dt	<=	188	;
						10'd19	:	dt	<=	188	;
						10'd20	:	dt	<=	187	;
						10'd21	:	dt	<=	186	;
						10'd22	:	dt	<=	184	;
						10'd23	:	dt	<=	184	;
						10'd24	:	dt	<=	182	;
						10'd25	:	dt	<=	182	;
						10'd26	:	dt	<=	181	;
						10'd27	:	dt	<=	180	;
						10'd28	:	dt	<=	193	;
						10'd29	:	dt	<=	194	;
						10'd30	:	dt	<=	195	;
						10'd31	:	dt	<=	195	;
						10'd32	:	dt	<=	195	;
						10'd33	:	dt	<=	195	;
						10'd34	:	dt	<=	195	;
						10'd35	:	dt	<=	195	;
						10'd36	:	dt	<=	195	;
						10'd37	:	dt	<=	194	;
						10'd38	:	dt	<=	194	;
						10'd39	:	dt	<=	195	;
						10'd40	:	dt	<=	196	;
						10'd41	:	dt	<=	194	;
						10'd42	:	dt	<=	193	;
						10'd43	:	dt	<=	193	;
						10'd44	:	dt	<=	193	;
						10'd45	:	dt	<=	195	;
						10'd46	:	dt	<=	192	;
						10'd47	:	dt	<=	189	;
						10'd48	:	dt	<=	188	;
						10'd49	:	dt	<=	187	;
						10'd50	:	dt	<=	187	;
						10'd51	:	dt	<=	186	;
						10'd52	:	dt	<=	185	;
						10'd53	:	dt	<=	184	;
						10'd54	:	dt	<=	183	;
						10'd55	:	dt	<=	181	;
						10'd56	:	dt	<=	198	;
						10'd57	:	dt	<=	197	;
						10'd58	:	dt	<=	198	;
						10'd59	:	dt	<=	197	;
						10'd60	:	dt	<=	197	;
						10'd61	:	dt	<=	198	;
						10'd62	:	dt	<=	197	;
						10'd63	:	dt	<=	197	;
						10'd64	:	dt	<=	197	;
						10'd65	:	dt	<=	198	;
						10'd66	:	dt	<=	197	;
						10'd67	:	dt	<=	195	;
						10'd68	:	dt	<=	193	;
						10'd69	:	dt	<=	199	;
						10'd70	:	dt	<=	198	;
						10'd71	:	dt	<=	189	;
						10'd72	:	dt	<=	164	;
						10'd73	:	dt	<=	155	;
						10'd74	:	dt	<=	190	;
						10'd75	:	dt	<=	195	;
						10'd76	:	dt	<=	194	;
						10'd77	:	dt	<=	193	;
						10'd78	:	dt	<=	188	;
						10'd79	:	dt	<=	188	;
						10'd80	:	dt	<=	188	;
						10'd81	:	dt	<=	187	;
						10'd82	:	dt	<=	186	;
						10'd83	:	dt	<=	185	;
						10'd84	:	dt	<=	200	;
						10'd85	:	dt	<=	199	;
						10'd86	:	dt	<=	199	;
						10'd87	:	dt	<=	200	;
						10'd88	:	dt	<=	199	;
						10'd89	:	dt	<=	199	;
						10'd90	:	dt	<=	199	;
						10'd91	:	dt	<=	199	;
						10'd92	:	dt	<=	199	;
						10'd93	:	dt	<=	198	;
						10'd94	:	dt	<=	197	;
						10'd95	:	dt	<=	183	;
						10'd96	:	dt	<=	159	;
						10'd97	:	dt	<=	161	;
						10'd98	:	dt	<=	197	;
						10'd99	:	dt	<=	192	;
						10'd100	:	dt	<=	163	;
						10'd101	:	dt	<=	122	;
						10'd102	:	dt	<=	145	;
						10'd103	:	dt	<=	193	;
						10'd104	:	dt	<=	159	;
						10'd105	:	dt	<=	168	;
						10'd106	:	dt	<=	193	;
						10'd107	:	dt	<=	190	;
						10'd108	:	dt	<=	189	;
						10'd109	:	dt	<=	189	;
						10'd110	:	dt	<=	187	;
						10'd111	:	dt	<=	186	;
						10'd112	:	dt	<=	202	;
						10'd113	:	dt	<=	201	;
						10'd114	:	dt	<=	201	;
						10'd115	:	dt	<=	202	;
						10'd116	:	dt	<=	202	;
						10'd117	:	dt	<=	201	;
						10'd118	:	dt	<=	201	;
						10'd119	:	dt	<=	201	;
						10'd120	:	dt	<=	201	;
						10'd121	:	dt	<=	200	;
						10'd122	:	dt	<=	204	;
						10'd123	:	dt	<=	207	;
						10'd124	:	dt	<=	182	;
						10'd125	:	dt	<=	152	;
						10'd126	:	dt	<=	141	;
						10'd127	:	dt	<=	187	;
						10'd128	:	dt	<=	181	;
						10'd129	:	dt	<=	145	;
						10'd130	:	dt	<=	108	;
						10'd131	:	dt	<=	159	;
						10'd132	:	dt	<=	152	;
						10'd133	:	dt	<=	111	;
						10'd134	:	dt	<=	157	;
						10'd135	:	dt	<=	200	;
						10'd136	:	dt	<=	189	;
						10'd137	:	dt	<=	191	;
						10'd138	:	dt	<=	189	;
						10'd139	:	dt	<=	188	;
						10'd140	:	dt	<=	202	;
						10'd141	:	dt	<=	202	;
						10'd142	:	dt	<=	203	;
						10'd143	:	dt	<=	204	;
						10'd144	:	dt	<=	204	;
						10'd145	:	dt	<=	203	;
						10'd146	:	dt	<=	203	;
						10'd147	:	dt	<=	204	;
						10'd148	:	dt	<=	202	;
						10'd149	:	dt	<=	196	;
						10'd150	:	dt	<=	193	;
						10'd151	:	dt	<=	196	;
						10'd152	:	dt	<=	203	;
						10'd153	:	dt	<=	181	;
						10'd154	:	dt	<=	136	;
						10'd155	:	dt	<=	136	;
						10'd156	:	dt	<=	186	;
						10'd157	:	dt	<=	163	;
						10'd158	:	dt	<=	110	;
						10'd159	:	dt	<=	136	;
						10'd160	:	dt	<=	162	;
						10'd161	:	dt	<=	116	;
						10'd162	:	dt	<=	107	;
						10'd163	:	dt	<=	198	;
						10'd164	:	dt	<=	192	;
						10'd165	:	dt	<=	193	;
						10'd166	:	dt	<=	191	;
						10'd167	:	dt	<=	190	;
						10'd168	:	dt	<=	205	;
						10'd169	:	dt	<=	204	;
						10'd170	:	dt	<=	204	;
						10'd171	:	dt	<=	205	;
						10'd172	:	dt	<=	205	;
						10'd173	:	dt	<=	206	;
						10'd174	:	dt	<=	205	;
						10'd175	:	dt	<=	207	;
						10'd176	:	dt	<=	198	;
						10'd177	:	dt	<=	187	;
						10'd178	:	dt	<=	185	;
						10'd179	:	dt	<=	143	;
						10'd180	:	dt	<=	163	;
						10'd181	:	dt	<=	180	;
						10'd182	:	dt	<=	123	;
						10'd183	:	dt	<=	105	;
						10'd184	:	dt	<=	183	;
						10'd185	:	dt	<=	162	;
						10'd186	:	dt	<=	110	;
						10'd187	:	dt	<=	117	;
						10'd188	:	dt	<=	164	;
						10'd189	:	dt	<=	131	;
						10'd190	:	dt	<=	95	;
						10'd191	:	dt	<=	193	;
						10'd192	:	dt	<=	195	;
						10'd193	:	dt	<=	193	;
						10'd194	:	dt	<=	192	;
						10'd195	:	dt	<=	191	;
						10'd196	:	dt	<=	206	;
						10'd197	:	dt	<=	206	;
						10'd198	:	dt	<=	207	;
						10'd199	:	dt	<=	207	;
						10'd200	:	dt	<=	207	;
						10'd201	:	dt	<=	206	;
						10'd202	:	dt	<=	207	;
						10'd203	:	dt	<=	206	;
						10'd204	:	dt	<=	201	;
						10'd205	:	dt	<=	198	;
						10'd206	:	dt	<=	189	;
						10'd207	:	dt	<=	142	;
						10'd208	:	dt	<=	120	;
						10'd209	:	dt	<=	161	;
						10'd210	:	dt	<=	115	;
						10'd211	:	dt	<=	99	;
						10'd212	:	dt	<=	164	;
						10'd213	:	dt	<=	133	;
						10'd214	:	dt	<=	90	;
						10'd215	:	dt	<=	137	;
						10'd216	:	dt	<=	169	;
						10'd217	:	dt	<=	137	;
						10'd218	:	dt	<=	107	;
						10'd219	:	dt	<=	200	;
						10'd220	:	dt	<=	197	;
						10'd221	:	dt	<=	196	;
						10'd222	:	dt	<=	195	;
						10'd223	:	dt	<=	195	;
						10'd224	:	dt	<=	207	;
						10'd225	:	dt	<=	207	;
						10'd226	:	dt	<=	208	;
						10'd227	:	dt	<=	207	;
						10'd228	:	dt	<=	208	;
						10'd229	:	dt	<=	208	;
						10'd230	:	dt	<=	208	;
						10'd231	:	dt	<=	209	;
						10'd232	:	dt	<=	194	;
						10'd233	:	dt	<=	154	;
						10'd234	:	dt	<=	181	;
						10'd235	:	dt	<=	158	;
						10'd236	:	dt	<=	114	;
						10'd237	:	dt	<=	141	;
						10'd238	:	dt	<=	146	;
						10'd239	:	dt	<=	97	;
						10'd240	:	dt	<=	133	;
						10'd241	:	dt	<=	120	;
						10'd242	:	dt	<=	78	;
						10'd243	:	dt	<=	144	;
						10'd244	:	dt	<=	143	;
						10'd245	:	dt	<=	102	;
						10'd246	:	dt	<=	123	;
						10'd247	:	dt	<=	209	;
						10'd248	:	dt	<=	197	;
						10'd249	:	dt	<=	198	;
						10'd250	:	dt	<=	198	;
						10'd251	:	dt	<=	196	;
						10'd252	:	dt	<=	209	;
						10'd253	:	dt	<=	208	;
						10'd254	:	dt	<=	209	;
						10'd255	:	dt	<=	209	;
						10'd256	:	dt	<=	209	;
						10'd257	:	dt	<=	209	;
						10'd258	:	dt	<=	209	;
						10'd259	:	dt	<=	208	;
						10'd260	:	dt	<=	207	;
						10'd261	:	dt	<=	154	;
						10'd262	:	dt	<=	140	;
						10'd263	:	dt	<=	182	;
						10'd264	:	dt	<=	144	;
						10'd265	:	dt	<=	124	;
						10'd266	:	dt	<=	172	;
						10'd267	:	dt	<=	105	;
						10'd268	:	dt	<=	112	;
						10'd269	:	dt	<=	137	;
						10'd270	:	dt	<=	133	;
						10'd271	:	dt	<=	138	;
						10'd272	:	dt	<=	105	;
						10'd273	:	dt	<=	68	;
						10'd274	:	dt	<=	145	;
						10'd275	:	dt	<=	212	;
						10'd276	:	dt	<=	199	;
						10'd277	:	dt	<=	200	;
						10'd278	:	dt	<=	199	;
						10'd279	:	dt	<=	198	;
						10'd280	:	dt	<=	210	;
						10'd281	:	dt	<=	210	;
						10'd282	:	dt	<=	209	;
						10'd283	:	dt	<=	210	;
						10'd284	:	dt	<=	211	;
						10'd285	:	dt	<=	209	;
						10'd286	:	dt	<=	208	;
						10'd287	:	dt	<=	211	;
						10'd288	:	dt	<=	196	;
						10'd289	:	dt	<=	138	;
						10'd290	:	dt	<=	113	;
						10'd291	:	dt	<=	172	;
						10'd292	:	dt	<=	148	;
						10'd293	:	dt	<=	164	;
						10'd294	:	dt	<=	171	;
						10'd295	:	dt	<=	151	;
						10'd296	:	dt	<=	154	;
						10'd297	:	dt	<=	153	;
						10'd298	:	dt	<=	179	;
						10'd299	:	dt	<=	150	;
						10'd300	:	dt	<=	94	;
						10'd301	:	dt	<=	72	;
						10'd302	:	dt	<=	182	;
						10'd303	:	dt	<=	207	;
						10'd304	:	dt	<=	201	;
						10'd305	:	dt	<=	202	;
						10'd306	:	dt	<=	200	;
						10'd307	:	dt	<=	199	;
						10'd308	:	dt	<=	210	;
						10'd309	:	dt	<=	210	;
						10'd310	:	dt	<=	211	;
						10'd311	:	dt	<=	211	;
						10'd312	:	dt	<=	210	;
						10'd313	:	dt	<=	210	;
						10'd314	:	dt	<=	210	;
						10'd315	:	dt	<=	212	;
						10'd316	:	dt	<=	196	;
						10'd317	:	dt	<=	171	;
						10'd318	:	dt	<=	168	;
						10'd319	:	dt	<=	140	;
						10'd320	:	dt	<=	94	;
						10'd321	:	dt	<=	181	;
						10'd322	:	dt	<=	171	;
						10'd323	:	dt	<=	160	;
						10'd324	:	dt	<=	169	;
						10'd325	:	dt	<=	157	;
						10'd326	:	dt	<=	167	;
						10'd327	:	dt	<=	141	;
						10'd328	:	dt	<=	102	;
						10'd329	:	dt	<=	95	;
						10'd330	:	dt	<=	206	;
						10'd331	:	dt	<=	204	;
						10'd332	:	dt	<=	203	;
						10'd333	:	dt	<=	203	;
						10'd334	:	dt	<=	202	;
						10'd335	:	dt	<=	200	;
						10'd336	:	dt	<=	211	;
						10'd337	:	dt	<=	211	;
						10'd338	:	dt	<=	211	;
						10'd339	:	dt	<=	211	;
						10'd340	:	dt	<=	212	;
						10'd341	:	dt	<=	212	;
						10'd342	:	dt	<=	211	;
						10'd343	:	dt	<=	211	;
						10'd344	:	dt	<=	207	;
						10'd345	:	dt	<=	193	;
						10'd346	:	dt	<=	156	;
						10'd347	:	dt	<=	120	;
						10'd348	:	dt	<=	88	;
						10'd349	:	dt	<=	117	;
						10'd350	:	dt	<=	148	;
						10'd351	:	dt	<=	137	;
						10'd352	:	dt	<=	140	;
						10'd353	:	dt	<=	137	;
						10'd354	:	dt	<=	131	;
						10'd355	:	dt	<=	130	;
						10'd356	:	dt	<=	120	;
						10'd357	:	dt	<=	93	;
						10'd358	:	dt	<=	179	;
						10'd359	:	dt	<=	213	;
						10'd360	:	dt	<=	204	;
						10'd361	:	dt	<=	204	;
						10'd362	:	dt	<=	203	;
						10'd363	:	dt	<=	201	;
						10'd364	:	dt	<=	212	;
						10'd365	:	dt	<=	212	;
						10'd366	:	dt	<=	212	;
						10'd367	:	dt	<=	212	;
						10'd368	:	dt	<=	213	;
						10'd369	:	dt	<=	212	;
						10'd370	:	dt	<=	211	;
						10'd371	:	dt	<=	210	;
						10'd372	:	dt	<=	208	;
						10'd373	:	dt	<=	181	;
						10'd374	:	dt	<=	142	;
						10'd375	:	dt	<=	109	;
						10'd376	:	dt	<=	99	;
						10'd377	:	dt	<=	97	;
						10'd378	:	dt	<=	115	;
						10'd379	:	dt	<=	125	;
						10'd380	:	dt	<=	125	;
						10'd381	:	dt	<=	120	;
						10'd382	:	dt	<=	112	;
						10'd383	:	dt	<=	141	;
						10'd384	:	dt	<=	135	;
						10'd385	:	dt	<=	108	;
						10'd386	:	dt	<=	110	;
						10'd387	:	dt	<=	211	;
						10'd388	:	dt	<=	206	;
						10'd389	:	dt	<=	205	;
						10'd390	:	dt	<=	205	;
						10'd391	:	dt	<=	204	;
						10'd392	:	dt	<=	213	;
						10'd393	:	dt	<=	213	;
						10'd394	:	dt	<=	213	;
						10'd395	:	dt	<=	213	;
						10'd396	:	dt	<=	213	;
						10'd397	:	dt	<=	214	;
						10'd398	:	dt	<=	212	;
						10'd399	:	dt	<=	210	;
						10'd400	:	dt	<=	200	;
						10'd401	:	dt	<=	164	;
						10'd402	:	dt	<=	130	;
						10'd403	:	dt	<=	106	;
						10'd404	:	dt	<=	103	;
						10'd405	:	dt	<=	122	;
						10'd406	:	dt	<=	127	;
						10'd407	:	dt	<=	155	;
						10'd408	:	dt	<=	164	;
						10'd409	:	dt	<=	159	;
						10'd410	:	dt	<=	141	;
						10'd411	:	dt	<=	148	;
						10'd412	:	dt	<=	149	;
						10'd413	:	dt	<=	140	;
						10'd414	:	dt	<=	92	;
						10'd415	:	dt	<=	160	;
						10'd416	:	dt	<=	217	;
						10'd417	:	dt	<=	203	;
						10'd418	:	dt	<=	205	;
						10'd419	:	dt	<=	204	;
						10'd420	:	dt	<=	214	;
						10'd421	:	dt	<=	215	;
						10'd422	:	dt	<=	215	;
						10'd423	:	dt	<=	215	;
						10'd424	:	dt	<=	215	;
						10'd425	:	dt	<=	215	;
						10'd426	:	dt	<=	213	;
						10'd427	:	dt	<=	207	;
						10'd428	:	dt	<=	201	;
						10'd429	:	dt	<=	175	;
						10'd430	:	dt	<=	143	;
						10'd431	:	dt	<=	113	;
						10'd432	:	dt	<=	115	;
						10'd433	:	dt	<=	122	;
						10'd434	:	dt	<=	146	;
						10'd435	:	dt	<=	183	;
						10'd436	:	dt	<=	183	;
						10'd437	:	dt	<=	197	;
						10'd438	:	dt	<=	184	;
						10'd439	:	dt	<=	159	;
						10'd440	:	dt	<=	186	;
						10'd441	:	dt	<=	161	;
						10'd442	:	dt	<=	109	;
						10'd443	:	dt	<=	106	;
						10'd444	:	dt	<=	214	;
						10'd445	:	dt	<=	206	;
						10'd446	:	dt	<=	206	;
						10'd447	:	dt	<=	205	;
						10'd448	:	dt	<=	216	;
						10'd449	:	dt	<=	216	;
						10'd450	:	dt	<=	215	;
						10'd451	:	dt	<=	216	;
						10'd452	:	dt	<=	216	;
						10'd453	:	dt	<=	216	;
						10'd454	:	dt	<=	215	;
						10'd455	:	dt	<=	205	;
						10'd456	:	dt	<=	202	;
						10'd457	:	dt	<=	178	;
						10'd458	:	dt	<=	144	;
						10'd459	:	dt	<=	111	;
						10'd460	:	dt	<=	111	;
						10'd461	:	dt	<=	131	;
						10'd462	:	dt	<=	164	;
						10'd463	:	dt	<=	193	;
						10'd464	:	dt	<=	194	;
						10'd465	:	dt	<=	205	;
						10'd466	:	dt	<=	209	;
						10'd467	:	dt	<=	191	;
						10'd468	:	dt	<=	175	;
						10'd469	:	dt	<=	160	;
						10'd470	:	dt	<=	106	;
						10'd471	:	dt	<=	101	;
						10'd472	:	dt	<=	213	;
						10'd473	:	dt	<=	208	;
						10'd474	:	dt	<=	207	;
						10'd475	:	dt	<=	206	;
						10'd476	:	dt	<=	216	;
						10'd477	:	dt	<=	217	;
						10'd478	:	dt	<=	216	;
						10'd479	:	dt	<=	216	;
						10'd480	:	dt	<=	216	;
						10'd481	:	dt	<=	217	;
						10'd482	:	dt	<=	216	;
						10'd483	:	dt	<=	199	;
						10'd484	:	dt	<=	200	;
						10'd485	:	dt	<=	188	;
						10'd486	:	dt	<=	152	;
						10'd487	:	dt	<=	119	;
						10'd488	:	dt	<=	117	;
						10'd489	:	dt	<=	133	;
						10'd490	:	dt	<=	167	;
						10'd491	:	dt	<=	201	;
						10'd492	:	dt	<=	202	;
						10'd493	:	dt	<=	210	;
						10'd494	:	dt	<=	200	;
						10'd495	:	dt	<=	185	;
						10'd496	:	dt	<=	165	;
						10'd497	:	dt	<=	134	;
						10'd498	:	dt	<=	88	;
						10'd499	:	dt	<=	134	;
						10'd500	:	dt	<=	221	;
						10'd501	:	dt	<=	207	;
						10'd502	:	dt	<=	208	;
						10'd503	:	dt	<=	207	;
						10'd504	:	dt	<=	216	;
						10'd505	:	dt	<=	216	;
						10'd506	:	dt	<=	217	;
						10'd507	:	dt	<=	217	;
						10'd508	:	dt	<=	217	;
						10'd509	:	dt	<=	217	;
						10'd510	:	dt	<=	217	;
						10'd511	:	dt	<=	195	;
						10'd512	:	dt	<=	199	;
						10'd513	:	dt	<=	195	;
						10'd514	:	dt	<=	159	;
						10'd515	:	dt	<=	132	;
						10'd516	:	dt	<=	126	;
						10'd517	:	dt	<=	129	;
						10'd518	:	dt	<=	176	;
						10'd519	:	dt	<=	207	;
						10'd520	:	dt	<=	211	;
						10'd521	:	dt	<=	210	;
						10'd522	:	dt	<=	192	;
						10'd523	:	dt	<=	173	;
						10'd524	:	dt	<=	155	;
						10'd525	:	dt	<=	118	;
						10'd526	:	dt	<=	80	;
						10'd527	:	dt	<=	183	;
						10'd528	:	dt	<=	218	;
						10'd529	:	dt	<=	209	;
						10'd530	:	dt	<=	209	;
						10'd531	:	dt	<=	208	;
						10'd532	:	dt	<=	217	;
						10'd533	:	dt	<=	217	;
						10'd534	:	dt	<=	218	;
						10'd535	:	dt	<=	218	;
						10'd536	:	dt	<=	218	;
						10'd537	:	dt	<=	218	;
						10'd538	:	dt	<=	220	;
						10'd539	:	dt	<=	195	;
						10'd540	:	dt	<=	193	;
						10'd541	:	dt	<=	196	;
						10'd542	:	dt	<=	169	;
						10'd543	:	dt	<=	139	;
						10'd544	:	dt	<=	128	;
						10'd545	:	dt	<=	134	;
						10'd546	:	dt	<=	183	;
						10'd547	:	dt	<=	212	;
						10'd548	:	dt	<=	211	;
						10'd549	:	dt	<=	202	;
						10'd550	:	dt	<=	184	;
						10'd551	:	dt	<=	164	;
						10'd552	:	dt	<=	147	;
						10'd553	:	dt	<=	100	;
						10'd554	:	dt	<=	101	;
						10'd555	:	dt	<=	217	;
						10'd556	:	dt	<=	211	;
						10'd557	:	dt	<=	211	;
						10'd558	:	dt	<=	210	;
						10'd559	:	dt	<=	209	;
						10'd560	:	dt	<=	217	;
						10'd561	:	dt	<=	217	;
						10'd562	:	dt	<=	218	;
						10'd563	:	dt	<=	219	;
						10'd564	:	dt	<=	218	;
						10'd565	:	dt	<=	218	;
						10'd566	:	dt	<=	221	;
						10'd567	:	dt	<=	199	;
						10'd568	:	dt	<=	180	;
						10'd569	:	dt	<=	187	;
						10'd570	:	dt	<=	169	;
						10'd571	:	dt	<=	142	;
						10'd572	:	dt	<=	129	;
						10'd573	:	dt	<=	140	;
						10'd574	:	dt	<=	192	;
						10'd575	:	dt	<=	209	;
						10'd576	:	dt	<=	200	;
						10'd577	:	dt	<=	193	;
						10'd578	:	dt	<=	174	;
						10'd579	:	dt	<=	150	;
						10'd580	:	dt	<=	134	;
						10'd581	:	dt	<=	85	;
						10'd582	:	dt	<=	150	;
						10'd583	:	dt	<=	224	;
						10'd584	:	dt	<=	209	;
						10'd585	:	dt	<=	212	;
						10'd586	:	dt	<=	210	;
						10'd587	:	dt	<=	210	;
						10'd588	:	dt	<=	217	;
						10'd589	:	dt	<=	217	;
						10'd590	:	dt	<=	217	;
						10'd591	:	dt	<=	218	;
						10'd592	:	dt	<=	218	;
						10'd593	:	dt	<=	218	;
						10'd594	:	dt	<=	221	;
						10'd595	:	dt	<=	212	;
						10'd596	:	dt	<=	177	;
						10'd597	:	dt	<=	187	;
						10'd598	:	dt	<=	175	;
						10'd599	:	dt	<=	145	;
						10'd600	:	dt	<=	139	;
						10'd601	:	dt	<=	145	;
						10'd602	:	dt	<=	196	;
						10'd603	:	dt	<=	200	;
						10'd604	:	dt	<=	191	;
						10'd605	:	dt	<=	182	;
						10'd606	:	dt	<=	161	;
						10'd607	:	dt	<=	137	;
						10'd608	:	dt	<=	113	;
						10'd609	:	dt	<=	85	;
						10'd610	:	dt	<=	201	;
						10'd611	:	dt	<=	219	;
						10'd612	:	dt	<=	213	;
						10'd613	:	dt	<=	212	;
						10'd614	:	dt	<=	211	;
						10'd615	:	dt	<=	211	;
						10'd616	:	dt	<=	216	;
						10'd617	:	dt	<=	216	;
						10'd618	:	dt	<=	217	;
						10'd619	:	dt	<=	218	;
						10'd620	:	dt	<=	217	;
						10'd621	:	dt	<=	217	;
						10'd622	:	dt	<=	217	;
						10'd623	:	dt	<=	220	;
						10'd624	:	dt	<=	189	;
						10'd625	:	dt	<=	185	;
						10'd626	:	dt	<=	180	;
						10'd627	:	dt	<=	159	;
						10'd628	:	dt	<=	157	;
						10'd629	:	dt	<=	142	;
						10'd630	:	dt	<=	192	;
						10'd631	:	dt	<=	191	;
						10'd632	:	dt	<=	188	;
						10'd633	:	dt	<=	168	;
						10'd634	:	dt	<=	146	;
						10'd635	:	dt	<=	127	;
						10'd636	:	dt	<=	87	;
						10'd637	:	dt	<=	125	;
						10'd638	:	dt	<=	225	;
						10'd639	:	dt	<=	212	;
						10'd640	:	dt	<=	214	;
						10'd641	:	dt	<=	212	;
						10'd642	:	dt	<=	210	;
						10'd643	:	dt	<=	210	;
						10'd644	:	dt	<=	216	;
						10'd645	:	dt	<=	216	;
						10'd646	:	dt	<=	217	;
						10'd647	:	dt	<=	218	;
						10'd648	:	dt	<=	217	;
						10'd649	:	dt	<=	217	;
						10'd650	:	dt	<=	217	;
						10'd651	:	dt	<=	222	;
						10'd652	:	dt	<=	204	;
						10'd653	:	dt	<=	181	;
						10'd654	:	dt	<=	181	;
						10'd655	:	dt	<=	171	;
						10'd656	:	dt	<=	157	;
						10'd657	:	dt	<=	133	;
						10'd658	:	dt	<=	174	;
						10'd659	:	dt	<=	182	;
						10'd660	:	dt	<=	179	;
						10'd661	:	dt	<=	156	;
						10'd662	:	dt	<=	128	;
						10'd663	:	dt	<=	106	;
						10'd664	:	dt	<=	79	;
						10'd665	:	dt	<=	194	;
						10'd666	:	dt	<=	218	;
						10'd667	:	dt	<=	211	;
						10'd668	:	dt	<=	211	;
						10'd669	:	dt	<=	211	;
						10'd670	:	dt	<=	210	;
						10'd671	:	dt	<=	210	;
						10'd672	:	dt	<=	217	;
						10'd673	:	dt	<=	216	;
						10'd674	:	dt	<=	218	;
						10'd675	:	dt	<=	218	;
						10'd676	:	dt	<=	218	;
						10'd677	:	dt	<=	218	;
						10'd678	:	dt	<=	218	;
						10'd679	:	dt	<=	221	;
						10'd680	:	dt	<=	211	;
						10'd681	:	dt	<=	186	;
						10'd682	:	dt	<=	178	;
						10'd683	:	dt	<=	165	;
						10'd684	:	dt	<=	151	;
						10'd685	:	dt	<=	135	;
						10'd686	:	dt	<=	156	;
						10'd687	:	dt	<=	164	;
						10'd688	:	dt	<=	153	;
						10'd689	:	dt	<=	130	;
						10'd690	:	dt	<=	107	;
						10'd691	:	dt	<=	73	;
						10'd692	:	dt	<=	141	;
						10'd693	:	dt	<=	226	;
						10'd694	:	dt	<=	212	;
						10'd695	:	dt	<=	214	;
						10'd696	:	dt	<=	213	;
						10'd697	:	dt	<=	212	;
						10'd698	:	dt	<=	211	;
						10'd699	:	dt	<=	210	;
						10'd700	:	dt	<=	217	;
						10'd701	:	dt	<=	218	;
						10'd702	:	dt	<=	218	;
						10'd703	:	dt	<=	218	;
						10'd704	:	dt	<=	218	;
						10'd705	:	dt	<=	218	;
						10'd706	:	dt	<=	219	;
						10'd707	:	dt	<=	221	;
						10'd708	:	dt	<=	213	;
						10'd709	:	dt	<=	193	;
						10'd710	:	dt	<=	181	;
						10'd711	:	dt	<=	163	;
						10'd712	:	dt	<=	148	;
						10'd713	:	dt	<=	137	;
						10'd714	:	dt	<=	145	;
						10'd715	:	dt	<=	154	;
						10'd716	:	dt	<=	133	;
						10'd717	:	dt	<=	108	;
						10'd718	:	dt	<=	84	;
						10'd719	:	dt	<=	89	;
						10'd720	:	dt	<=	213	;
						10'd721	:	dt	<=	218	;
						10'd722	:	dt	<=	216	;
						10'd723	:	dt	<=	215	;
						10'd724	:	dt	<=	213	;
						10'd725	:	dt	<=	212	;
						10'd726	:	dt	<=	211	;
						10'd727	:	dt	<=	210	;
						10'd728	:	dt	<=	217	;
						10'd729	:	dt	<=	219	;
						10'd730	:	dt	<=	219	;
						10'd731	:	dt	<=	219	;
						10'd732	:	dt	<=	218	;
						10'd733	:	dt	<=	218	;
						10'd734	:	dt	<=	220	;
						10'd735	:	dt	<=	222	;
						10'd736	:	dt	<=	203	;
						10'd737	:	dt	<=	194	;
						10'd738	:	dt	<=	182	;
						10'd739	:	dt	<=	167	;
						10'd740	:	dt	<=	155	;
						10'd741	:	dt	<=	148	;
						10'd742	:	dt	<=	143	;
						10'd743	:	dt	<=	149	;
						10'd744	:	dt	<=	136	;
						10'd745	:	dt	<=	106	;
						10'd746	:	dt	<=	72	;
						10'd747	:	dt	<=	150	;
						10'd748	:	dt	<=	229	;
						10'd749	:	dt	<=	214	;
						10'd750	:	dt	<=	217	;
						10'd751	:	dt	<=	215	;
						10'd752	:	dt	<=	213	;
						10'd753	:	dt	<=	212	;
						10'd754	:	dt	<=	211	;
						10'd755	:	dt	<=	212	;
						10'd756	:	dt	<=	217	;
						10'd757	:	dt	<=	217	;
						10'd758	:	dt	<=	218	;
						10'd759	:	dt	<=	218	;
						10'd760	:	dt	<=	219	;
						10'd761	:	dt	<=	218	;
						10'd762	:	dt	<=	220	;
						10'd763	:	dt	<=	218	;
						10'd764	:	dt	<=	190	;
						10'd765	:	dt	<=	193	;
						10'd766	:	dt	<=	185	;
						10'd767	:	dt	<=	178	;
						10'd768	:	dt	<=	175	;
						10'd769	:	dt	<=	162	;
						10'd770	:	dt	<=	150	;
						10'd771	:	dt	<=	142	;
						10'd772	:	dt	<=	128	;
						10'd773	:	dt	<=	97	;
						10'd774	:	dt	<=	81	;
						10'd775	:	dt	<=	192	;
						10'd776	:	dt	<=	223	;
						10'd777	:	dt	<=	216	;
						10'd778	:	dt	<=	216	;
						10'd779	:	dt	<=	215	;
						10'd780	:	dt	<=	214	;
						10'd781	:	dt	<=	213	;
						10'd782	:	dt	<=	212	;
						10'd783	:	dt	<=	204	;
					endcase
				end
				5'd5	:	begin
					case (cnt)
						10'd0	:	dt	<=	126	;
						10'd1	:	dt	<=	128	;
						10'd2	:	dt	<=	131	;
						10'd3	:	dt	<=	132	;
						10'd4	:	dt	<=	133	;
						10'd5	:	dt	<=	134	;
						10'd6	:	dt	<=	135	;
						10'd7	:	dt	<=	135	;
						10'd8	:	dt	<=	136	;
						10'd9	:	dt	<=	138	;
						10'd10	:	dt	<=	137	;
						10'd11	:	dt	<=	137	;
						10'd12	:	dt	<=	138	;
						10'd13	:	dt	<=	138	;
						10'd14	:	dt	<=	139	;
						10'd15	:	dt	<=	137	;
						10'd16	:	dt	<=	142	;
						10'd17	:	dt	<=	140	;
						10'd18	:	dt	<=	138	;
						10'd19	:	dt	<=	139	;
						10'd20	:	dt	<=	137	;
						10'd21	:	dt	<=	137	;
						10'd22	:	dt	<=	136	;
						10'd23	:	dt	<=	135	;
						10'd24	:	dt	<=	134	;
						10'd25	:	dt	<=	133	;
						10'd26	:	dt	<=	134	;
						10'd27	:	dt	<=	132	;
						10'd28	:	dt	<=	129	;
						10'd29	:	dt	<=	132	;
						10'd30	:	dt	<=	134	;
						10'd31	:	dt	<=	135	;
						10'd32	:	dt	<=	135	;
						10'd33	:	dt	<=	137	;
						10'd34	:	dt	<=	139	;
						10'd35	:	dt	<=	139	;
						10'd36	:	dt	<=	139	;
						10'd37	:	dt	<=	140	;
						10'd38	:	dt	<=	141	;
						10'd39	:	dt	<=	141	;
						10'd40	:	dt	<=	142	;
						10'd41	:	dt	<=	143	;
						10'd42	:	dt	<=	142	;
						10'd43	:	dt	<=	142	;
						10'd44	:	dt	<=	116	;
						10'd45	:	dt	<=	138	;
						10'd46	:	dt	<=	141	;
						10'd47	:	dt	<=	140	;
						10'd48	:	dt	<=	141	;
						10'd49	:	dt	<=	140	;
						10'd50	:	dt	<=	139	;
						10'd51	:	dt	<=	138	;
						10'd52	:	dt	<=	137	;
						10'd53	:	dt	<=	136	;
						10'd54	:	dt	<=	136	;
						10'd55	:	dt	<=	134	;
						10'd56	:	dt	<=	133	;
						10'd57	:	dt	<=	135	;
						10'd58	:	dt	<=	138	;
						10'd59	:	dt	<=	139	;
						10'd60	:	dt	<=	139	;
						10'd61	:	dt	<=	141	;
						10'd62	:	dt	<=	142	;
						10'd63	:	dt	<=	143	;
						10'd64	:	dt	<=	142	;
						10'd65	:	dt	<=	143	;
						10'd66	:	dt	<=	145	;
						10'd67	:	dt	<=	145	;
						10'd68	:	dt	<=	143	;
						10'd69	:	dt	<=	145	;
						10'd70	:	dt	<=	145	;
						10'd71	:	dt	<=	158	;
						10'd72	:	dt	<=	94	;
						10'd73	:	dt	<=	118	;
						10'd74	:	dt	<=	151	;
						10'd75	:	dt	<=	143	;
						10'd76	:	dt	<=	144	;
						10'd77	:	dt	<=	144	;
						10'd78	:	dt	<=	142	;
						10'd79	:	dt	<=	141	;
						10'd80	:	dt	<=	141	;
						10'd81	:	dt	<=	140	;
						10'd82	:	dt	<=	139	;
						10'd83	:	dt	<=	138	;
						10'd84	:	dt	<=	137	;
						10'd85	:	dt	<=	139	;
						10'd86	:	dt	<=	142	;
						10'd87	:	dt	<=	142	;
						10'd88	:	dt	<=	142	;
						10'd89	:	dt	<=	144	;
						10'd90	:	dt	<=	146	;
						10'd91	:	dt	<=	146	;
						10'd92	:	dt	<=	146	;
						10'd93	:	dt	<=	147	;
						10'd94	:	dt	<=	147	;
						10'd95	:	dt	<=	147	;
						10'd96	:	dt	<=	148	;
						10'd97	:	dt	<=	117	;
						10'd98	:	dt	<=	128	;
						10'd99	:	dt	<=	168	;
						10'd100	:	dt	<=	101	;
						10'd101	:	dt	<=	98	;
						10'd102	:	dt	<=	157	;
						10'd103	:	dt	<=	146	;
						10'd104	:	dt	<=	147	;
						10'd105	:	dt	<=	146	;
						10'd106	:	dt	<=	146	;
						10'd107	:	dt	<=	145	;
						10'd108	:	dt	<=	144	;
						10'd109	:	dt	<=	143	;
						10'd110	:	dt	<=	142	;
						10'd111	:	dt	<=	141	;
						10'd112	:	dt	<=	140	;
						10'd113	:	dt	<=	142	;
						10'd114	:	dt	<=	145	;
						10'd115	:	dt	<=	146	;
						10'd116	:	dt	<=	147	;
						10'd117	:	dt	<=	148	;
						10'd118	:	dt	<=	149	;
						10'd119	:	dt	<=	149	;
						10'd120	:	dt	<=	149	;
						10'd121	:	dt	<=	151	;
						10'd122	:	dt	<=	151	;
						10'd123	:	dt	<=	149	;
						10'd124	:	dt	<=	161	;
						10'd125	:	dt	<=	114	;
						10'd126	:	dt	<=	99	;
						10'd127	:	dt	<=	174	;
						10'd128	:	dt	<=	99	;
						10'd129	:	dt	<=	84	;
						10'd130	:	dt	<=	162	;
						10'd131	:	dt	<=	149	;
						10'd132	:	dt	<=	151	;
						10'd133	:	dt	<=	149	;
						10'd134	:	dt	<=	148	;
						10'd135	:	dt	<=	147	;
						10'd136	:	dt	<=	146	;
						10'd137	:	dt	<=	146	;
						10'd138	:	dt	<=	145	;
						10'd139	:	dt	<=	144	;
						10'd140	:	dt	<=	143	;
						10'd141	:	dt	<=	145	;
						10'd142	:	dt	<=	149	;
						10'd143	:	dt	<=	150	;
						10'd144	:	dt	<=	150	;
						10'd145	:	dt	<=	151	;
						10'd146	:	dt	<=	153	;
						10'd147	:	dt	<=	153	;
						10'd148	:	dt	<=	154	;
						10'd149	:	dt	<=	153	;
						10'd150	:	dt	<=	154	;
						10'd151	:	dt	<=	152	;
						10'd152	:	dt	<=	167	;
						10'd153	:	dt	<=	126	;
						10'd154	:	dt	<=	88	;
						10'd155	:	dt	<=	169	;
						10'd156	:	dt	<=	99	;
						10'd157	:	dt	<=	87	;
						10'd158	:	dt	<=	164	;
						10'd159	:	dt	<=	152	;
						10'd160	:	dt	<=	153	;
						10'd161	:	dt	<=	152	;
						10'd162	:	dt	<=	151	;
						10'd163	:	dt	<=	150	;
						10'd164	:	dt	<=	149	;
						10'd165	:	dt	<=	148	;
						10'd166	:	dt	<=	148	;
						10'd167	:	dt	<=	147	;
						10'd168	:	dt	<=	145	;
						10'd169	:	dt	<=	147	;
						10'd170	:	dt	<=	151	;
						10'd171	:	dt	<=	152	;
						10'd172	:	dt	<=	153	;
						10'd173	:	dt	<=	155	;
						10'd174	:	dt	<=	155	;
						10'd175	:	dt	<=	155	;
						10'd176	:	dt	<=	151	;
						10'd177	:	dt	<=	154	;
						10'd178	:	dt	<=	158	;
						10'd179	:	dt	<=	155	;
						10'd180	:	dt	<=	170	;
						10'd181	:	dt	<=	130	;
						10'd182	:	dt	<=	79	;
						10'd183	:	dt	<=	166	;
						10'd184	:	dt	<=	111	;
						10'd185	:	dt	<=	93	;
						10'd186	:	dt	<=	166	;
						10'd187	:	dt	<=	156	;
						10'd188	:	dt	<=	157	;
						10'd189	:	dt	<=	156	;
						10'd190	:	dt	<=	155	;
						10'd191	:	dt	<=	153	;
						10'd192	:	dt	<=	152	;
						10'd193	:	dt	<=	152	;
						10'd194	:	dt	<=	152	;
						10'd195	:	dt	<=	150	;
						10'd196	:	dt	<=	149	;
						10'd197	:	dt	<=	150	;
						10'd198	:	dt	<=	153	;
						10'd199	:	dt	<=	155	;
						10'd200	:	dt	<=	155	;
						10'd201	:	dt	<=	158	;
						10'd202	:	dt	<=	157	;
						10'd203	:	dt	<=	163	;
						10'd204	:	dt	<=	129	;
						10'd205	:	dt	<=	120	;
						10'd206	:	dt	<=	166	;
						10'd207	:	dt	<=	156	;
						10'd208	:	dt	<=	171	;
						10'd209	:	dt	<=	140	;
						10'd210	:	dt	<=	82	;
						10'd211	:	dt	<=	162	;
						10'd212	:	dt	<=	102	;
						10'd213	:	dt	<=	97	;
						10'd214	:	dt	<=	168	;
						10'd215	:	dt	<=	158	;
						10'd216	:	dt	<=	160	;
						10'd217	:	dt	<=	158	;
						10'd218	:	dt	<=	162	;
						10'd219	:	dt	<=	160	;
						10'd220	:	dt	<=	154	;
						10'd221	:	dt	<=	154	;
						10'd222	:	dt	<=	154	;
						10'd223	:	dt	<=	152	;
						10'd224	:	dt	<=	151	;
						10'd225	:	dt	<=	152	;
						10'd226	:	dt	<=	156	;
						10'd227	:	dt	<=	158	;
						10'd228	:	dt	<=	159	;
						10'd229	:	dt	<=	159	;
						10'd230	:	dt	<=	158	;
						10'd231	:	dt	<=	164	;
						10'd232	:	dt	<=	139	;
						10'd233	:	dt	<=	91	;
						10'd234	:	dt	<=	165	;
						10'd235	:	dt	<=	159	;
						10'd236	:	dt	<=	174	;
						10'd237	:	dt	<=	144	;
						10'd238	:	dt	<=	71	;
						10'd239	:	dt	<=	156	;
						10'd240	:	dt	<=	96	;
						10'd241	:	dt	<=	100	;
						10'd242	:	dt	<=	171	;
						10'd243	:	dt	<=	161	;
						10'd244	:	dt	<=	161	;
						10'd245	:	dt	<=	158	;
						10'd246	:	dt	<=	128	;
						10'd247	:	dt	<=	145	;
						10'd248	:	dt	<=	162	;
						10'd249	:	dt	<=	156	;
						10'd250	:	dt	<=	155	;
						10'd251	:	dt	<=	155	;
						10'd252	:	dt	<=	152	;
						10'd253	:	dt	<=	155	;
						10'd254	:	dt	<=	159	;
						10'd255	:	dt	<=	160	;
						10'd256	:	dt	<=	161	;
						10'd257	:	dt	<=	161	;
						10'd258	:	dt	<=	160	;
						10'd259	:	dt	<=	168	;
						10'd260	:	dt	<=	158	;
						10'd261	:	dt	<=	76	;
						10'd262	:	dt	<=	159	;
						10'd263	:	dt	<=	164	;
						10'd264	:	dt	<=	172	;
						10'd265	:	dt	<=	142	;
						10'd266	:	dt	<=	63	;
						10'd267	:	dt	<=	155	;
						10'd268	:	dt	<=	117	;
						10'd269	:	dt	<=	100	;
						10'd270	:	dt	<=	174	;
						10'd271	:	dt	<=	159	;
						10'd272	:	dt	<=	164	;
						10'd273	:	dt	<=	164	;
						10'd274	:	dt	<=	126	;
						10'd275	:	dt	<=	103	;
						10'd276	:	dt	<=	162	;
						10'd277	:	dt	<=	161	;
						10'd278	:	dt	<=	158	;
						10'd279	:	dt	<=	157	;
						10'd280	:	dt	<=	153	;
						10'd281	:	dt	<=	157	;
						10'd282	:	dt	<=	160	;
						10'd283	:	dt	<=	162	;
						10'd284	:	dt	<=	162	;
						10'd285	:	dt	<=	162	;
						10'd286	:	dt	<=	164	;
						10'd287	:	dt	<=	167	;
						10'd288	:	dt	<=	158	;
						10'd289	:	dt	<=	78	;
						10'd290	:	dt	<=	158	;
						10'd291	:	dt	<=	167	;
						10'd292	:	dt	<=	167	;
						10'd293	:	dt	<=	156	;
						10'd294	:	dt	<=	73	;
						10'd295	:	dt	<=	133	;
						10'd296	:	dt	<=	129	;
						10'd297	:	dt	<=	102	;
						10'd298	:	dt	<=	172	;
						10'd299	:	dt	<=	157	;
						10'd300	:	dt	<=	148	;
						10'd301	:	dt	<=	130	;
						10'd302	:	dt	<=	156	;
						10'd303	:	dt	<=	132	;
						10'd304	:	dt	<=	129	;
						10'd305	:	dt	<=	163	;
						10'd306	:	dt	<=	161	;
						10'd307	:	dt	<=	159	;
						10'd308	:	dt	<=	157	;
						10'd309	:	dt	<=	159	;
						10'd310	:	dt	<=	162	;
						10'd311	:	dt	<=	164	;
						10'd312	:	dt	<=	164	;
						10'd313	:	dt	<=	165	;
						10'd314	:	dt	<=	166	;
						10'd315	:	dt	<=	167	;
						10'd316	:	dt	<=	173	;
						10'd317	:	dt	<=	89	;
						10'd318	:	dt	<=	139	;
						10'd319	:	dt	<=	172	;
						10'd320	:	dt	<=	162	;
						10'd321	:	dt	<=	163	;
						10'd322	:	dt	<=	79	;
						10'd323	:	dt	<=	98	;
						10'd324	:	dt	<=	132	;
						10'd325	:	dt	<=	111	;
						10'd326	:	dt	<=	170	;
						10'd327	:	dt	<=	160	;
						10'd328	:	dt	<=	142	;
						10'd329	:	dt	<=	54	;
						10'd330	:	dt	<=	125	;
						10'd331	:	dt	<=	150	;
						10'd332	:	dt	<=	102	;
						10'd333	:	dt	<=	150	;
						10'd334	:	dt	<=	167	;
						10'd335	:	dt	<=	162	;
						10'd336	:	dt	<=	159	;
						10'd337	:	dt	<=	161	;
						10'd338	:	dt	<=	166	;
						10'd339	:	dt	<=	165	;
						10'd340	:	dt	<=	167	;
						10'd341	:	dt	<=	167	;
						10'd342	:	dt	<=	167	;
						10'd343	:	dt	<=	168	;
						10'd344	:	dt	<=	178	;
						10'd345	:	dt	<=	118	;
						10'd346	:	dt	<=	112	;
						10'd347	:	dt	<=	175	;
						10'd348	:	dt	<=	164	;
						10'd349	:	dt	<=	167	;
						10'd350	:	dt	<=	82	;
						10'd351	:	dt	<=	91	;
						10'd352	:	dt	<=	129	;
						10'd353	:	dt	<=	110	;
						10'd354	:	dt	<=	160	;
						10'd355	:	dt	<=	156	;
						10'd356	:	dt	<=	130	;
						10'd357	:	dt	<=	96	;
						10'd358	:	dt	<=	157	;
						10'd359	:	dt	<=	130	;
						10'd360	:	dt	<=	106	;
						10'd361	:	dt	<=	169	;
						10'd362	:	dt	<=	165	;
						10'd363	:	dt	<=	164	;
						10'd364	:	dt	<=	159	;
						10'd365	:	dt	<=	162	;
						10'd366	:	dt	<=	166	;
						10'd367	:	dt	<=	167	;
						10'd368	:	dt	<=	168	;
						10'd369	:	dt	<=	168	;
						10'd370	:	dt	<=	170	;
						10'd371	:	dt	<=	169	;
						10'd372	:	dt	<=	164	;
						10'd373	:	dt	<=	168	;
						10'd374	:	dt	<=	132	;
						10'd375	:	dt	<=	141	;
						10'd376	:	dt	<=	162	;
						10'd377	:	dt	<=	153	;
						10'd378	:	dt	<=	103	;
						10'd379	:	dt	<=	113	;
						10'd380	:	dt	<=	117	;
						10'd381	:	dt	<=	96	;
						10'd382	:	dt	<=	133	;
						10'd383	:	dt	<=	143	;
						10'd384	:	dt	<=	107	;
						10'd385	:	dt	<=	147	;
						10'd386	:	dt	<=	172	;
						10'd387	:	dt	<=	99	;
						10'd388	:	dt	<=	139	;
						10'd389	:	dt	<=	174	;
						10'd390	:	dt	<=	165	;
						10'd391	:	dt	<=	166	;
						10'd392	:	dt	<=	161	;
						10'd393	:	dt	<=	164	;
						10'd394	:	dt	<=	167	;
						10'd395	:	dt	<=	170	;
						10'd396	:	dt	<=	171	;
						10'd397	:	dt	<=	171	;
						10'd398	:	dt	<=	170	;
						10'd399	:	dt	<=	173	;
						10'd400	:	dt	<=	160	;
						10'd401	:	dt	<=	173	;
						10'd402	:	dt	<=	162	;
						10'd403	:	dt	<=	129	;
						10'd404	:	dt	<=	132	;
						10'd405	:	dt	<=	132	;
						10'd406	:	dt	<=	109	;
						10'd407	:	dt	<=	109	;
						10'd408	:	dt	<=	108	;
						10'd409	:	dt	<=	99	;
						10'd410	:	dt	<=	135	;
						10'd411	:	dt	<=	142	;
						10'd412	:	dt	<=	111	;
						10'd413	:	dt	<=	163	;
						10'd414	:	dt	<=	154	;
						10'd415	:	dt	<=	77	;
						10'd416	:	dt	<=	156	;
						10'd417	:	dt	<=	172	;
						10'd418	:	dt	<=	167	;
						10'd419	:	dt	<=	167	;
						10'd420	:	dt	<=	165	;
						10'd421	:	dt	<=	167	;
						10'd422	:	dt	<=	168	;
						10'd423	:	dt	<=	171	;
						10'd424	:	dt	<=	172	;
						10'd425	:	dt	<=	173	;
						10'd426	:	dt	<=	173	;
						10'd427	:	dt	<=	174	;
						10'd428	:	dt	<=	169	;
						10'd429	:	dt	<=	170	;
						10'd430	:	dt	<=	182	;
						10'd431	:	dt	<=	150	;
						10'd432	:	dt	<=	125	;
						10'd433	:	dt	<=	124	;
						10'd434	:	dt	<=	100	;
						10'd435	:	dt	<=	106	;
						10'd436	:	dt	<=	103	;
						10'd437	:	dt	<=	102	;
						10'd438	:	dt	<=	130	;
						10'd439	:	dt	<=	138	;
						10'd440	:	dt	<=	124	;
						10'd441	:	dt	<=	178	;
						10'd442	:	dt	<=	130	;
						10'd443	:	dt	<=	64	;
						10'd444	:	dt	<=	168	;
						10'd445	:	dt	<=	172	;
						10'd446	:	dt	<=	170	;
						10'd447	:	dt	<=	169	;
						10'd448	:	dt	<=	165	;
						10'd449	:	dt	<=	168	;
						10'd450	:	dt	<=	170	;
						10'd451	:	dt	<=	171	;
						10'd452	:	dt	<=	172	;
						10'd453	:	dt	<=	174	;
						10'd454	:	dt	<=	175	;
						10'd455	:	dt	<=	174	;
						10'd456	:	dt	<=	175	;
						10'd457	:	dt	<=	172	;
						10'd458	:	dt	<=	195	;
						10'd459	:	dt	<=	170	;
						10'd460	:	dt	<=	114	;
						10'd461	:	dt	<=	110	;
						10'd462	:	dt	<=	94	;
						10'd463	:	dt	<=	89	;
						10'd464	:	dt	<=	98	;
						10'd465	:	dt	<=	105	;
						10'd466	:	dt	<=	127	;
						10'd467	:	dt	<=	134	;
						10'd468	:	dt	<=	124	;
						10'd469	:	dt	<=	182	;
						10'd470	:	dt	<=	126	;
						10'd471	:	dt	<=	80	;
						10'd472	:	dt	<=	180	;
						10'd473	:	dt	<=	171	;
						10'd474	:	dt	<=	171	;
						10'd475	:	dt	<=	171	;
						10'd476	:	dt	<=	166	;
						10'd477	:	dt	<=	169	;
						10'd478	:	dt	<=	171	;
						10'd479	:	dt	<=	172	;
						10'd480	:	dt	<=	173	;
						10'd481	:	dt	<=	174	;
						10'd482	:	dt	<=	175	;
						10'd483	:	dt	<=	176	;
						10'd484	:	dt	<=	177	;
						10'd485	:	dt	<=	174	;
						10'd486	:	dt	<=	197	;
						10'd487	:	dt	<=	179	;
						10'd488	:	dt	<=	119	;
						10'd489	:	dt	<=	86	;
						10'd490	:	dt	<=	87	;
						10'd491	:	dt	<=	81	;
						10'd492	:	dt	<=	94	;
						10'd493	:	dt	<=	118	;
						10'd494	:	dt	<=	136	;
						10'd495	:	dt	<=	123	;
						10'd496	:	dt	<=	116	;
						10'd497	:	dt	<=	177	;
						10'd498	:	dt	<=	127	;
						10'd499	:	dt	<=	94	;
						10'd500	:	dt	<=	183	;
						10'd501	:	dt	<=	172	;
						10'd502	:	dt	<=	173	;
						10'd503	:	dt	<=	173	;
						10'd504	:	dt	<=	169	;
						10'd505	:	dt	<=	172	;
						10'd506	:	dt	<=	172	;
						10'd507	:	dt	<=	174	;
						10'd508	:	dt	<=	175	;
						10'd509	:	dt	<=	174	;
						10'd510	:	dt	<=	177	;
						10'd511	:	dt	<=	178	;
						10'd512	:	dt	<=	178	;
						10'd513	:	dt	<=	175	;
						10'd514	:	dt	<=	192	;
						10'd515	:	dt	<=	176	;
						10'd516	:	dt	<=	126	;
						10'd517	:	dt	<=	87	;
						10'd518	:	dt	<=	86	;
						10'd519	:	dt	<=	82	;
						10'd520	:	dt	<=	109	;
						10'd521	:	dt	<=	130	;
						10'd522	:	dt	<=	147	;
						10'd523	:	dt	<=	159	;
						10'd524	:	dt	<=	128	;
						10'd525	:	dt	<=	164	;
						10'd526	:	dt	<=	128	;
						10'd527	:	dt	<=	100	;
						10'd528	:	dt	<=	184	;
						10'd529	:	dt	<=	174	;
						10'd530	:	dt	<=	173	;
						10'd531	:	dt	<=	173	;
						10'd532	:	dt	<=	169	;
						10'd533	:	dt	<=	172	;
						10'd534	:	dt	<=	173	;
						10'd535	:	dt	<=	173	;
						10'd536	:	dt	<=	176	;
						10'd537	:	dt	<=	178	;
						10'd538	:	dt	<=	179	;
						10'd539	:	dt	<=	178	;
						10'd540	:	dt	<=	181	;
						10'd541	:	dt	<=	175	;
						10'd542	:	dt	<=	189	;
						10'd543	:	dt	<=	171	;
						10'd544	:	dt	<=	126	;
						10'd545	:	dt	<=	89	;
						10'd546	:	dt	<=	80	;
						10'd547	:	dt	<=	90	;
						10'd548	:	dt	<=	121	;
						10'd549	:	dt	<=	137	;
						10'd550	:	dt	<=	164	;
						10'd551	:	dt	<=	175	;
						10'd552	:	dt	<=	141	;
						10'd553	:	dt	<=	140	;
						10'd554	:	dt	<=	108	;
						10'd555	:	dt	<=	95	;
						10'd556	:	dt	<=	184	;
						10'd557	:	dt	<=	176	;
						10'd558	:	dt	<=	175	;
						10'd559	:	dt	<=	173	;
						10'd560	:	dt	<=	171	;
						10'd561	:	dt	<=	173	;
						10'd562	:	dt	<=	174	;
						10'd563	:	dt	<=	175	;
						10'd564	:	dt	<=	177	;
						10'd565	:	dt	<=	179	;
						10'd566	:	dt	<=	179	;
						10'd567	:	dt	<=	179	;
						10'd568	:	dt	<=	181	;
						10'd569	:	dt	<=	174	;
						10'd570	:	dt	<=	189	;
						10'd571	:	dt	<=	171	;
						10'd572	:	dt	<=	134	;
						10'd573	:	dt	<=	91	;
						10'd574	:	dt	<=	80	;
						10'd575	:	dt	<=	98	;
						10'd576	:	dt	<=	134	;
						10'd577	:	dt	<=	159	;
						10'd578	:	dt	<=	164	;
						10'd579	:	dt	<=	167	;
						10'd580	:	dt	<=	153	;
						10'd581	:	dt	<=	114	;
						10'd582	:	dt	<=	73	;
						10'd583	:	dt	<=	82	;
						10'd584	:	dt	<=	185	;
						10'd585	:	dt	<=	176	;
						10'd586	:	dt	<=	177	;
						10'd587	:	dt	<=	177	;
						10'd588	:	dt	<=	172	;
						10'd589	:	dt	<=	173	;
						10'd590	:	dt	<=	174	;
						10'd591	:	dt	<=	177	;
						10'd592	:	dt	<=	178	;
						10'd593	:	dt	<=	179	;
						10'd594	:	dt	<=	180	;
						10'd595	:	dt	<=	180	;
						10'd596	:	dt	<=	183	;
						10'd597	:	dt	<=	174	;
						10'd598	:	dt	<=	186	;
						10'd599	:	dt	<=	172	;
						10'd600	:	dt	<=	138	;
						10'd601	:	dt	<=	93	;
						10'd602	:	dt	<=	82	;
						10'd603	:	dt	<=	97	;
						10'd604	:	dt	<=	143	;
						10'd605	:	dt	<=	172	;
						10'd606	:	dt	<=	169	;
						10'd607	:	dt	<=	160	;
						10'd608	:	dt	<=	132	;
						10'd609	:	dt	<=	89	;
						10'd610	:	dt	<=	44	;
						10'd611	:	dt	<=	108	;
						10'd612	:	dt	<=	189	;
						10'd613	:	dt	<=	176	;
						10'd614	:	dt	<=	178	;
						10'd615	:	dt	<=	178	;
						10'd616	:	dt	<=	171	;
						10'd617	:	dt	<=	173	;
						10'd618	:	dt	<=	177	;
						10'd619	:	dt	<=	178	;
						10'd620	:	dt	<=	179	;
						10'd621	:	dt	<=	180	;
						10'd622	:	dt	<=	181	;
						10'd623	:	dt	<=	182	;
						10'd624	:	dt	<=	185	;
						10'd625	:	dt	<=	178	;
						10'd626	:	dt	<=	179	;
						10'd627	:	dt	<=	170	;
						10'd628	:	dt	<=	137	;
						10'd629	:	dt	<=	95	;
						10'd630	:	dt	<=	88	;
						10'd631	:	dt	<=	90	;
						10'd632	:	dt	<=	152	;
						10'd633	:	dt	<=	180	;
						10'd634	:	dt	<=	167	;
						10'd635	:	dt	<=	141	;
						10'd636	:	dt	<=	112	;
						10'd637	:	dt	<=	65	;
						10'd638	:	dt	<=	64	;
						10'd639	:	dt	<=	176	;
						10'd640	:	dt	<=	183	;
						10'd641	:	dt	<=	179	;
						10'd642	:	dt	<=	179	;
						10'd643	:	dt	<=	178	;
						10'd644	:	dt	<=	173	;
						10'd645	:	dt	<=	174	;
						10'd646	:	dt	<=	178	;
						10'd647	:	dt	<=	179	;
						10'd648	:	dt	<=	179	;
						10'd649	:	dt	<=	180	;
						10'd650	:	dt	<=	182	;
						10'd651	:	dt	<=	183	;
						10'd652	:	dt	<=	186	;
						10'd653	:	dt	<=	175	;
						10'd654	:	dt	<=	165	;
						10'd655	:	dt	<=	168	;
						10'd656	:	dt	<=	137	;
						10'd657	:	dt	<=	100	;
						10'd658	:	dt	<=	96	;
						10'd659	:	dt	<=	88	;
						10'd660	:	dt	<=	149	;
						10'd661	:	dt	<=	168	;
						10'd662	:	dt	<=	147	;
						10'd663	:	dt	<=	122	;
						10'd664	:	dt	<=	92	;
						10'd665	:	dt	<=	50	;
						10'd666	:	dt	<=	144	;
						10'd667	:	dt	<=	193	;
						10'd668	:	dt	<=	181	;
						10'd669	:	dt	<=	181	;
						10'd670	:	dt	<=	180	;
						10'd671	:	dt	<=	179	;
						10'd672	:	dt	<=	173	;
						10'd673	:	dt	<=	174	;
						10'd674	:	dt	<=	177	;
						10'd675	:	dt	<=	179	;
						10'd676	:	dt	<=	180	;
						10'd677	:	dt	<=	180	;
						10'd678	:	dt	<=	183	;
						10'd679	:	dt	<=	182	;
						10'd680	:	dt	<=	187	;
						10'd681	:	dt	<=	177	;
						10'd682	:	dt	<=	158	;
						10'd683	:	dt	<=	161	;
						10'd684	:	dt	<=	130	;
						10'd685	:	dt	<=	111	;
						10'd686	:	dt	<=	101	;
						10'd687	:	dt	<=	91	;
						10'd688	:	dt	<=	136	;
						10'd689	:	dt	<=	150	;
						10'd690	:	dt	<=	135	;
						10'd691	:	dt	<=	112	;
						10'd692	:	dt	<=	62	;
						10'd693	:	dt	<=	87	;
						10'd694	:	dt	<=	192	;
						10'd695	:	dt	<=	183	;
						10'd696	:	dt	<=	185	;
						10'd697	:	dt	<=	183	;
						10'd698	:	dt	<=	181	;
						10'd699	:	dt	<=	180	;
						10'd700	:	dt	<=	173	;
						10'd701	:	dt	<=	174	;
						10'd702	:	dt	<=	177	;
						10'd703	:	dt	<=	178	;
						10'd704	:	dt	<=	179	;
						10'd705	:	dt	<=	179	;
						10'd706	:	dt	<=	181	;
						10'd707	:	dt	<=	182	;
						10'd708	:	dt	<=	184	;
						10'd709	:	dt	<=	179	;
						10'd710	:	dt	<=	156	;
						10'd711	:	dt	<=	151	;
						10'd712	:	dt	<=	124	;
						10'd713	:	dt	<=	116	;
						10'd714	:	dt	<=	96	;
						10'd715	:	dt	<=	88	;
						10'd716	:	dt	<=	128	;
						10'd717	:	dt	<=	138	;
						10'd718	:	dt	<=	126	;
						10'd719	:	dt	<=	81	;
						10'd720	:	dt	<=	49	;
						10'd721	:	dt	<=	164	;
						10'd722	:	dt	<=	190	;
						10'd723	:	dt	<=	184	;
						10'd724	:	dt	<=	185	;
						10'd725	:	dt	<=	184	;
						10'd726	:	dt	<=	182	;
						10'd727	:	dt	<=	181	;
						10'd728	:	dt	<=	172	;
						10'd729	:	dt	<=	174	;
						10'd730	:	dt	<=	177	;
						10'd731	:	dt	<=	178	;
						10'd732	:	dt	<=	178	;
						10'd733	:	dt	<=	178	;
						10'd734	:	dt	<=	180	;
						10'd735	:	dt	<=	182	;
						10'd736	:	dt	<=	184	;
						10'd737	:	dt	<=	177	;
						10'd738	:	dt	<=	160	;
						10'd739	:	dt	<=	154	;
						10'd740	:	dt	<=	128	;
						10'd741	:	dt	<=	114	;
						10'd742	:	dt	<=	97	;
						10'd743	:	dt	<=	78	;
						10'd744	:	dt	<=	114	;
						10'd745	:	dt	<=	112	;
						10'd746	:	dt	<=	89	;
						10'd747	:	dt	<=	48	;
						10'd748	:	dt	<=	133	;
						10'd749	:	dt	<=	194	;
						10'd750	:	dt	<=	182	;
						10'd751	:	dt	<=	185	;
						10'd752	:	dt	<=	184	;
						10'd753	:	dt	<=	184	;
						10'd754	:	dt	<=	182	;
						10'd755	:	dt	<=	181	;
						10'd756	:	dt	<=	172	;
						10'd757	:	dt	<=	174	;
						10'd758	:	dt	<=	177	;
						10'd759	:	dt	<=	178	;
						10'd760	:	dt	<=	178	;
						10'd761	:	dt	<=	179	;
						10'd762	:	dt	<=	181	;
						10'd763	:	dt	<=	183	;
						10'd764	:	dt	<=	187	;
						10'd765	:	dt	<=	175	;
						10'd766	:	dt	<=	165	;
						10'd767	:	dt	<=	154	;
						10'd768	:	dt	<=	118	;
						10'd769	:	dt	<=	107	;
						10'd770	:	dt	<=	100	;
						10'd771	:	dt	<=	75	;
						10'd772	:	dt	<=	96	;
						10'd773	:	dt	<=	83	;
						10'd774	:	dt	<=	47	;
						10'd775	:	dt	<=	104	;
						10'd776	:	dt	<=	194	;
						10'd777	:	dt	<=	183	;
						10'd778	:	dt	<=	186	;
						10'd779	:	dt	<=	184	;
						10'd780	:	dt	<=	184	;
						10'd781	:	dt	<=	184	;
						10'd782	:	dt	<=	182	;
						10'd783	:	dt	<=	180	;
					endcase
				end
				5'd6	:	begin
					case (cnt)
						10'd0	:	dt	<=	149	;
						10'd1	:	dt	<=	149	;
						10'd2	:	dt	<=	150	;
						10'd3	:	dt	<=	150	;
						10'd4	:	dt	<=	150	;
						10'd5	:	dt	<=	151	;
						10'd6	:	dt	<=	151	;
						10'd7	:	dt	<=	150	;
						10'd8	:	dt	<=	151	;
						10'd9	:	dt	<=	152	;
						10'd10	:	dt	<=	152	;
						10'd11	:	dt	<=	152	;
						10'd12	:	dt	<=	152	;
						10'd13	:	dt	<=	152	;
						10'd14	:	dt	<=	153	;
						10'd15	:	dt	<=	153	;
						10'd16	:	dt	<=	151	;
						10'd17	:	dt	<=	152	;
						10'd18	:	dt	<=	152	;
						10'd19	:	dt	<=	153	;
						10'd20	:	dt	<=	152	;
						10'd21	:	dt	<=	152	;
						10'd22	:	dt	<=	151	;
						10'd23	:	dt	<=	151	;
						10'd24	:	dt	<=	150	;
						10'd25	:	dt	<=	150	;
						10'd26	:	dt	<=	150	;
						10'd27	:	dt	<=	149	;
						10'd28	:	dt	<=	150	;
						10'd29	:	dt	<=	150	;
						10'd30	:	dt	<=	150	;
						10'd31	:	dt	<=	152	;
						10'd32	:	dt	<=	152	;
						10'd33	:	dt	<=	151	;
						10'd34	:	dt	<=	152	;
						10'd35	:	dt	<=	152	;
						10'd36	:	dt	<=	152	;
						10'd37	:	dt	<=	152	;
						10'd38	:	dt	<=	152	;
						10'd39	:	dt	<=	153	;
						10'd40	:	dt	<=	154	;
						10'd41	:	dt	<=	153	;
						10'd42	:	dt	<=	154	;
						10'd43	:	dt	<=	154	;
						10'd44	:	dt	<=	153	;
						10'd45	:	dt	<=	154	;
						10'd46	:	dt	<=	153	;
						10'd47	:	dt	<=	154	;
						10'd48	:	dt	<=	153	;
						10'd49	:	dt	<=	153	;
						10'd50	:	dt	<=	152	;
						10'd51	:	dt	<=	152	;
						10'd52	:	dt	<=	152	;
						10'd53	:	dt	<=	151	;
						10'd54	:	dt	<=	150	;
						10'd55	:	dt	<=	151	;
						10'd56	:	dt	<=	150	;
						10'd57	:	dt	<=	151	;
						10'd58	:	dt	<=	151	;
						10'd59	:	dt	<=	152	;
						10'd60	:	dt	<=	152	;
						10'd61	:	dt	<=	152	;
						10'd62	:	dt	<=	153	;
						10'd63	:	dt	<=	153	;
						10'd64	:	dt	<=	152	;
						10'd65	:	dt	<=	152	;
						10'd66	:	dt	<=	152	;
						10'd67	:	dt	<=	153	;
						10'd68	:	dt	<=	154	;
						10'd69	:	dt	<=	154	;
						10'd70	:	dt	<=	155	;
						10'd71	:	dt	<=	155	;
						10'd72	:	dt	<=	154	;
						10'd73	:	dt	<=	154	;
						10'd74	:	dt	<=	155	;
						10'd75	:	dt	<=	155	;
						10'd76	:	dt	<=	155	;
						10'd77	:	dt	<=	155	;
						10'd78	:	dt	<=	154	;
						10'd79	:	dt	<=	153	;
						10'd80	:	dt	<=	153	;
						10'd81	:	dt	<=	151	;
						10'd82	:	dt	<=	151	;
						10'd83	:	dt	<=	152	;
						10'd84	:	dt	<=	150	;
						10'd85	:	dt	<=	151	;
						10'd86	:	dt	<=	151	;
						10'd87	:	dt	<=	152	;
						10'd88	:	dt	<=	152	;
						10'd89	:	dt	<=	152	;
						10'd90	:	dt	<=	154	;
						10'd91	:	dt	<=	154	;
						10'd92	:	dt	<=	154	;
						10'd93	:	dt	<=	154	;
						10'd94	:	dt	<=	154	;
						10'd95	:	dt	<=	153	;
						10'd96	:	dt	<=	154	;
						10'd97	:	dt	<=	155	;
						10'd98	:	dt	<=	156	;
						10'd99	:	dt	<=	157	;
						10'd100	:	dt	<=	157	;
						10'd101	:	dt	<=	156	;
						10'd102	:	dt	<=	155	;
						10'd103	:	dt	<=	156	;
						10'd104	:	dt	<=	155	;
						10'd105	:	dt	<=	154	;
						10'd106	:	dt	<=	154	;
						10'd107	:	dt	<=	155	;
						10'd108	:	dt	<=	152	;
						10'd109	:	dt	<=	154	;
						10'd110	:	dt	<=	153	;
						10'd111	:	dt	<=	153	;
						10'd112	:	dt	<=	151	;
						10'd113	:	dt	<=	152	;
						10'd114	:	dt	<=	152	;
						10'd115	:	dt	<=	152	;
						10'd116	:	dt	<=	154	;
						10'd117	:	dt	<=	154	;
						10'd118	:	dt	<=	154	;
						10'd119	:	dt	<=	154	;
						10'd120	:	dt	<=	154	;
						10'd121	:	dt	<=	155	;
						10'd122	:	dt	<=	157	;
						10'd123	:	dt	<=	156	;
						10'd124	:	dt	<=	156	;
						10'd125	:	dt	<=	156	;
						10'd126	:	dt	<=	154	;
						10'd127	:	dt	<=	150	;
						10'd128	:	dt	<=	146	;
						10'd129	:	dt	<=	147	;
						10'd130	:	dt	<=	146	;
						10'd131	:	dt	<=	147	;
						10'd132	:	dt	<=	143	;
						10'd133	:	dt	<=	137	;
						10'd134	:	dt	<=	126	;
						10'd135	:	dt	<=	126	;
						10'd136	:	dt	<=	142	;
						10'd137	:	dt	<=	139	;
						10'd138	:	dt	<=	152	;
						10'd139	:	dt	<=	154	;
						10'd140	:	dt	<=	152	;
						10'd141	:	dt	<=	153	;
						10'd142	:	dt	<=	153	;
						10'd143	:	dt	<=	154	;
						10'd144	:	dt	<=	154	;
						10'd145	:	dt	<=	155	;
						10'd146	:	dt	<=	154	;
						10'd147	:	dt	<=	155	;
						10'd148	:	dt	<=	155	;
						10'd149	:	dt	<=	154	;
						10'd150	:	dt	<=	153	;
						10'd151	:	dt	<=	150	;
						10'd152	:	dt	<=	144	;
						10'd153	:	dt	<=	143	;
						10'd154	:	dt	<=	145	;
						10'd155	:	dt	<=	139	;
						10'd156	:	dt	<=	142	;
						10'd157	:	dt	<=	144	;
						10'd158	:	dt	<=	157	;
						10'd159	:	dt	<=	157	;
						10'd160	:	dt	<=	147	;
						10'd161	:	dt	<=	139	;
						10'd162	:	dt	<=	128	;
						10'd163	:	dt	<=	119	;
						10'd164	:	dt	<=	130	;
						10'd165	:	dt	<=	113	;
						10'd166	:	dt	<=	147	;
						10'd167	:	dt	<=	156	;
						10'd168	:	dt	<=	151	;
						10'd169	:	dt	<=	153	;
						10'd170	:	dt	<=	153	;
						10'd171	:	dt	<=	155	;
						10'd172	:	dt	<=	155	;
						10'd173	:	dt	<=	156	;
						10'd174	:	dt	<=	155	;
						10'd175	:	dt	<=	152	;
						10'd176	:	dt	<=	145	;
						10'd177	:	dt	<=	139	;
						10'd178	:	dt	<=	141	;
						10'd179	:	dt	<=	141	;
						10'd180	:	dt	<=	141	;
						10'd181	:	dt	<=	153	;
						10'd182	:	dt	<=	153	;
						10'd183	:	dt	<=	143	;
						10'd184	:	dt	<=	135	;
						10'd185	:	dt	<=	137	;
						10'd186	:	dt	<=	139	;
						10'd187	:	dt	<=	133	;
						10'd188	:	dt	<=	121	;
						10'd189	:	dt	<=	107	;
						10'd190	:	dt	<=	101	;
						10'd191	:	dt	<=	104	;
						10'd192	:	dt	<=	110	;
						10'd193	:	dt	<=	127	;
						10'd194	:	dt	<=	157	;
						10'd195	:	dt	<=	156	;
						10'd196	:	dt	<=	151	;
						10'd197	:	dt	<=	152	;
						10'd198	:	dt	<=	153	;
						10'd199	:	dt	<=	155	;
						10'd200	:	dt	<=	155	;
						10'd201	:	dt	<=	154	;
						10'd202	:	dt	<=	151	;
						10'd203	:	dt	<=	146	;
						10'd204	:	dt	<=	139	;
						10'd205	:	dt	<=	131	;
						10'd206	:	dt	<=	130	;
						10'd207	:	dt	<=	134	;
						10'd208	:	dt	<=	137	;
						10'd209	:	dt	<=	132	;
						10'd210	:	dt	<=	125	;
						10'd211	:	dt	<=	111	;
						10'd212	:	dt	<=	101	;
						10'd213	:	dt	<=	94	;
						10'd214	:	dt	<=	95	;
						10'd215	:	dt	<=	105	;
						10'd216	:	dt	<=	113	;
						10'd217	:	dt	<=	122	;
						10'd218	:	dt	<=	133	;
						10'd219	:	dt	<=	145	;
						10'd220	:	dt	<=	153	;
						10'd221	:	dt	<=	157	;
						10'd222	:	dt	<=	156	;
						10'd223	:	dt	<=	156	;
						10'd224	:	dt	<=	152	;
						10'd225	:	dt	<=	152	;
						10'd226	:	dt	<=	154	;
						10'd227	:	dt	<=	152	;
						10'd228	:	dt	<=	151	;
						10'd229	:	dt	<=	150	;
						10'd230	:	dt	<=	149	;
						10'd231	:	dt	<=	149	;
						10'd232	:	dt	<=	139	;
						10'd233	:	dt	<=	122	;
						10'd234	:	dt	<=	104	;
						10'd235	:	dt	<=	98	;
						10'd236	:	dt	<=	92	;
						10'd237	:	dt	<=	82	;
						10'd238	:	dt	<=	81	;
						10'd239	:	dt	<=	81	;
						10'd240	:	dt	<=	85	;
						10'd241	:	dt	<=	114	;
						10'd242	:	dt	<=	145	;
						10'd243	:	dt	<=	157	;
						10'd244	:	dt	<=	160	;
						10'd245	:	dt	<=	162	;
						10'd246	:	dt	<=	161	;
						10'd247	:	dt	<=	159	;
						10'd248	:	dt	<=	157	;
						10'd249	:	dt	<=	156	;
						10'd250	:	dt	<=	156	;
						10'd251	:	dt	<=	156	;
						10'd252	:	dt	<=	151	;
						10'd253	:	dt	<=	151	;
						10'd254	:	dt	<=	150	;
						10'd255	:	dt	<=	146	;
						10'd256	:	dt	<=	145	;
						10'd257	:	dt	<=	147	;
						10'd258	:	dt	<=	148	;
						10'd259	:	dt	<=	147	;
						10'd260	:	dt	<=	145	;
						10'd261	:	dt	<=	132	;
						10'd262	:	dt	<=	97	;
						10'd263	:	dt	<=	71	;
						10'd264	:	dt	<=	62	;
						10'd265	:	dt	<=	66	;
						10'd266	:	dt	<=	88	;
						10'd267	:	dt	<=	116	;
						10'd268	:	dt	<=	145	;
						10'd269	:	dt	<=	162	;
						10'd270	:	dt	<=	160	;
						10'd271	:	dt	<=	159	;
						10'd272	:	dt	<=	157	;
						10'd273	:	dt	<=	155	;
						10'd274	:	dt	<=	156	;
						10'd275	:	dt	<=	157	;
						10'd276	:	dt	<=	157	;
						10'd277	:	dt	<=	156	;
						10'd278	:	dt	<=	155	;
						10'd279	:	dt	<=	155	;
						10'd280	:	dt	<=	151	;
						10'd281	:	dt	<=	145	;
						10'd282	:	dt	<=	144	;
						10'd283	:	dt	<=	145	;
						10'd284	:	dt	<=	147	;
						10'd285	:	dt	<=	145	;
						10'd286	:	dt	<=	147	;
						10'd287	:	dt	<=	150	;
						10'd288	:	dt	<=	150	;
						10'd289	:	dt	<=	124	;
						10'd290	:	dt	<=	92	;
						10'd291	:	dt	<=	68	;
						10'd292	:	dt	<=	63	;
						10'd293	:	dt	<=	67	;
						10'd294	:	dt	<=	86	;
						10'd295	:	dt	<=	159	;
						10'd296	:	dt	<=	163	;
						10'd297	:	dt	<=	155	;
						10'd298	:	dt	<=	158	;
						10'd299	:	dt	<=	157	;
						10'd300	:	dt	<=	156	;
						10'd301	:	dt	<=	156	;
						10'd302	:	dt	<=	157	;
						10'd303	:	dt	<=	156	;
						10'd304	:	dt	<=	156	;
						10'd305	:	dt	<=	156	;
						10'd306	:	dt	<=	155	;
						10'd307	:	dt	<=	154	;
						10'd308	:	dt	<=	143	;
						10'd309	:	dt	<=	144	;
						10'd310	:	dt	<=	145	;
						10'd311	:	dt	<=	145	;
						10'd312	:	dt	<=	143	;
						10'd313	:	dt	<=	147	;
						10'd314	:	dt	<=	152	;
						10'd315	:	dt	<=	152	;
						10'd316	:	dt	<=	128	;
						10'd317	:	dt	<=	90	;
						10'd318	:	dt	<=	79	;
						10'd319	:	dt	<=	68	;
						10'd320	:	dt	<=	64	;
						10'd321	:	dt	<=	70	;
						10'd322	:	dt	<=	67	;
						10'd323	:	dt	<=	84	;
						10'd324	:	dt	<=	147	;
						10'd325	:	dt	<=	164	;
						10'd326	:	dt	<=	157	;
						10'd327	:	dt	<=	158	;
						10'd328	:	dt	<=	157	;
						10'd329	:	dt	<=	157	;
						10'd330	:	dt	<=	157	;
						10'd331	:	dt	<=	156	;
						10'd332	:	dt	<=	157	;
						10'd333	:	dt	<=	156	;
						10'd334	:	dt	<=	156	;
						10'd335	:	dt	<=	155	;
						10'd336	:	dt	<=	145	;
						10'd337	:	dt	<=	146	;
						10'd338	:	dt	<=	143	;
						10'd339	:	dt	<=	145	;
						10'd340	:	dt	<=	145	;
						10'd341	:	dt	<=	150	;
						10'd342	:	dt	<=	149	;
						10'd343	:	dt	<=	149	;
						10'd344	:	dt	<=	139	;
						10'd345	:	dt	<=	118	;
						10'd346	:	dt	<=	85	;
						10'd347	:	dt	<=	62	;
						10'd348	:	dt	<=	62	;
						10'd349	:	dt	<=	75	;
						10'd350	:	dt	<=	73	;
						10'd351	:	dt	<=	62	;
						10'd352	:	dt	<=	67	;
						10'd353	:	dt	<=	140	;
						10'd354	:	dt	<=	164	;
						10'd355	:	dt	<=	157	;
						10'd356	:	dt	<=	158	;
						10'd357	:	dt	<=	158	;
						10'd358	:	dt	<=	158	;
						10'd359	:	dt	<=	158	;
						10'd360	:	dt	<=	157	;
						10'd361	:	dt	<=	157	;
						10'd362	:	dt	<=	156	;
						10'd363	:	dt	<=	156	;
						10'd364	:	dt	<=	150	;
						10'd365	:	dt	<=	147	;
						10'd366	:	dt	<=	144	;
						10'd367	:	dt	<=	147	;
						10'd368	:	dt	<=	149	;
						10'd369	:	dt	<=	148	;
						10'd370	:	dt	<=	149	;
						10'd371	:	dt	<=	158	;
						10'd372	:	dt	<=	158	;
						10'd373	:	dt	<=	136	;
						10'd374	:	dt	<=	94	;
						10'd375	:	dt	<=	63	;
						10'd376	:	dt	<=	58	;
						10'd377	:	dt	<=	69	;
						10'd378	:	dt	<=	85	;
						10'd379	:	dt	<=	82	;
						10'd380	:	dt	<=	67	;
						10'd381	:	dt	<=	70	;
						10'd382	:	dt	<=	156	;
						10'd383	:	dt	<=	160	;
						10'd384	:	dt	<=	159	;
						10'd385	:	dt	<=	160	;
						10'd386	:	dt	<=	159	;
						10'd387	:	dt	<=	158	;
						10'd388	:	dt	<=	157	;
						10'd389	:	dt	<=	156	;
						10'd390	:	dt	<=	156	;
						10'd391	:	dt	<=	156	;
						10'd392	:	dt	<=	147	;
						10'd393	:	dt	<=	148	;
						10'd394	:	dt	<=	147	;
						10'd395	:	dt	<=	145	;
						10'd396	:	dt	<=	148	;
						10'd397	:	dt	<=	152	;
						10'd398	:	dt	<=	151	;
						10'd399	:	dt	<=	160	;
						10'd400	:	dt	<=	153	;
						10'd401	:	dt	<=	119	;
						10'd402	:	dt	<=	86	;
						10'd403	:	dt	<=	66	;
						10'd404	:	dt	<=	64	;
						10'd405	:	dt	<=	63	;
						10'd406	:	dt	<=	69	;
						10'd407	:	dt	<=	75	;
						10'd408	:	dt	<=	78	;
						10'd409	:	dt	<=	57	;
						10'd410	:	dt	<=	130	;
						10'd411	:	dt	<=	165	;
						10'd412	:	dt	<=	158	;
						10'd413	:	dt	<=	159	;
						10'd414	:	dt	<=	158	;
						10'd415	:	dt	<=	159	;
						10'd416	:	dt	<=	158	;
						10'd417	:	dt	<=	157	;
						10'd418	:	dt	<=	157	;
						10'd419	:	dt	<=	157	;
						10'd420	:	dt	<=	149	;
						10'd421	:	dt	<=	148	;
						10'd422	:	dt	<=	146	;
						10'd423	:	dt	<=	145	;
						10'd424	:	dt	<=	147	;
						10'd425	:	dt	<=	149	;
						10'd426	:	dt	<=	146	;
						10'd427	:	dt	<=	151	;
						10'd428	:	dt	<=	144	;
						10'd429	:	dt	<=	110	;
						10'd430	:	dt	<=	78	;
						10'd431	:	dt	<=	65	;
						10'd432	:	dt	<=	66	;
						10'd433	:	dt	<=	66	;
						10'd434	:	dt	<=	58	;
						10'd435	:	dt	<=	59	;
						10'd436	:	dt	<=	64	;
						10'd437	:	dt	<=	79	;
						10'd438	:	dt	<=	150	;
						10'd439	:	dt	<=	165	;
						10'd440	:	dt	<=	162	;
						10'd441	:	dt	<=	162	;
						10'd442	:	dt	<=	162	;
						10'd443	:	dt	<=	162	;
						10'd444	:	dt	<=	161	;
						10'd445	:	dt	<=	161	;
						10'd446	:	dt	<=	158	;
						10'd447	:	dt	<=	156	;
						10'd448	:	dt	<=	151	;
						10'd449	:	dt	<=	146	;
						10'd450	:	dt	<=	143	;
						10'd451	:	dt	<=	141	;
						10'd452	:	dt	<=	138	;
						10'd453	:	dt	<=	140	;
						10'd454	:	dt	<=	142	;
						10'd455	:	dt	<=	146	;
						10'd456	:	dt	<=	144	;
						10'd457	:	dt	<=	121	;
						10'd458	:	dt	<=	84	;
						10'd459	:	dt	<=	56	;
						10'd460	:	dt	<=	62	;
						10'd461	:	dt	<=	70	;
						10'd462	:	dt	<=	71	;
						10'd463	:	dt	<=	68	;
						10'd464	:	dt	<=	57	;
						10'd465	:	dt	<=	117	;
						10'd466	:	dt	<=	144	;
						10'd467	:	dt	<=	144	;
						10'd468	:	dt	<=	147	;
						10'd469	:	dt	<=	149	;
						10'd470	:	dt	<=	152	;
						10'd471	:	dt	<=	150	;
						10'd472	:	dt	<=	146	;
						10'd473	:	dt	<=	146	;
						10'd474	:	dt	<=	154	;
						10'd475	:	dt	<=	160	;
						10'd476	:	dt	<=	147	;
						10'd477	:	dt	<=	144	;
						10'd478	:	dt	<=	143	;
						10'd479	:	dt	<=	142	;
						10'd480	:	dt	<=	140	;
						10'd481	:	dt	<=	142	;
						10'd482	:	dt	<=	146	;
						10'd483	:	dt	<=	151	;
						10'd484	:	dt	<=	154	;
						10'd485	:	dt	<=	131	;
						10'd486	:	dt	<=	85	;
						10'd487	:	dt	<=	59	;
						10'd488	:	dt	<=	51	;
						10'd489	:	dt	<=	60	;
						10'd490	:	dt	<=	85	;
						10'd491	:	dt	<=	69	;
						10'd492	:	dt	<=	64	;
						10'd493	:	dt	<=	76	;
						10'd494	:	dt	<=	75	;
						10'd495	:	dt	<=	79	;
						10'd496	:	dt	<=	81	;
						10'd497	:	dt	<=	79	;
						10'd498	:	dt	<=	76	;
						10'd499	:	dt	<=	83	;
						10'd500	:	dt	<=	112	;
						10'd501	:	dt	<=	141	;
						10'd502	:	dt	<=	163	;
						10'd503	:	dt	<=	163	;
						10'd504	:	dt	<=	144	;
						10'd505	:	dt	<=	148	;
						10'd506	:	dt	<=	147	;
						10'd507	:	dt	<=	145	;
						10'd508	:	dt	<=	145	;
						10'd509	:	dt	<=	148	;
						10'd510	:	dt	<=	150	;
						10'd511	:	dt	<=	155	;
						10'd512	:	dt	<=	151	;
						10'd513	:	dt	<=	119	;
						10'd514	:	dt	<=	74	;
						10'd515	:	dt	<=	62	;
						10'd516	:	dt	<=	63	;
						10'd517	:	dt	<=	55	;
						10'd518	:	dt	<=	62	;
						10'd519	:	dt	<=	72	;
						10'd520	:	dt	<=	73	;
						10'd521	:	dt	<=	77	;
						10'd522	:	dt	<=	74	;
						10'd523	:	dt	<=	73	;
						10'd524	:	dt	<=	68	;
						10'd525	:	dt	<=	88	;
						10'd526	:	dt	<=	113	;
						10'd527	:	dt	<=	138	;
						10'd528	:	dt	<=	162	;
						10'd529	:	dt	<=	162	;
						10'd530	:	dt	<=	168	;
						10'd531	:	dt	<=	168	;
						10'd532	:	dt	<=	146	;
						10'd533	:	dt	<=	146	;
						10'd534	:	dt	<=	142	;
						10'd535	:	dt	<=	141	;
						10'd536	:	dt	<=	141	;
						10'd537	:	dt	<=	138	;
						10'd538	:	dt	<=	134	;
						10'd539	:	dt	<=	142	;
						10'd540	:	dt	<=	124	;
						10'd541	:	dt	<=	96	;
						10'd542	:	dt	<=	75	;
						10'd543	:	dt	<=	67	;
						10'd544	:	dt	<=	65	;
						10'd545	:	dt	<=	63	;
						10'd546	:	dt	<=	62	;
						10'd547	:	dt	<=	78	;
						10'd548	:	dt	<=	87	;
						10'd549	:	dt	<=	76	;
						10'd550	:	dt	<=	84	;
						10'd551	:	dt	<=	96	;
						10'd552	:	dt	<=	126	;
						10'd553	:	dt	<=	162	;
						10'd554	:	dt	<=	172	;
						10'd555	:	dt	<=	155	;
						10'd556	:	dt	<=	144	;
						10'd557	:	dt	<=	149	;
						10'd558	:	dt	<=	151	;
						10'd559	:	dt	<=	161	;
						10'd560	:	dt	<=	142	;
						10'd561	:	dt	<=	136	;
						10'd562	:	dt	<=	132	;
						10'd563	:	dt	<=	134	;
						10'd564	:	dt	<=	127	;
						10'd565	:	dt	<=	119	;
						10'd566	:	dt	<=	118	;
						10'd567	:	dt	<=	119	;
						10'd568	:	dt	<=	103	;
						10'd569	:	dt	<=	87	;
						10'd570	:	dt	<=	77	;
						10'd571	:	dt	<=	73	;
						10'd572	:	dt	<=	70	;
						10'd573	:	dt	<=	62	;
						10'd574	:	dt	<=	64	;
						10'd575	:	dt	<=	72	;
						10'd576	:	dt	<=	93	;
						10'd577	:	dt	<=	134	;
						10'd578	:	dt	<=	155	;
						10'd579	:	dt	<=	160	;
						10'd580	:	dt	<=	166	;
						10'd581	:	dt	<=	156	;
						10'd582	:	dt	<=	150	;
						10'd583	:	dt	<=	151	;
						10'd584	:	dt	<=	143	;
						10'd585	:	dt	<=	136	;
						10'd586	:	dt	<=	145	;
						10'd587	:	dt	<=	149	;
						10'd588	:	dt	<=	130	;
						10'd589	:	dt	<=	132	;
						10'd590	:	dt	<=	127	;
						10'd591	:	dt	<=	120	;
						10'd592	:	dt	<=	114	;
						10'd593	:	dt	<=	110	;
						10'd594	:	dt	<=	109	;
						10'd595	:	dt	<=	105	;
						10'd596	:	dt	<=	91	;
						10'd597	:	dt	<=	77	;
						10'd598	:	dt	<=	74	;
						10'd599	:	dt	<=	75	;
						10'd600	:	dt	<=	74	;
						10'd601	:	dt	<=	65	;
						10'd602	:	dt	<=	73	;
						10'd603	:	dt	<=	113	;
						10'd604	:	dt	<=	166	;
						10'd605	:	dt	<=	177	;
						10'd606	:	dt	<=	170	;
						10'd607	:	dt	<=	161	;
						10'd608	:	dt	<=	152	;
						10'd609	:	dt	<=	141	;
						10'd610	:	dt	<=	134	;
						10'd611	:	dt	<=	136	;
						10'd612	:	dt	<=	140	;
						10'd613	:	dt	<=	133	;
						10'd614	:	dt	<=	127	;
						10'd615	:	dt	<=	130	;
						10'd616	:	dt	<=	113	;
						10'd617	:	dt	<=	116	;
						10'd618	:	dt	<=	115	;
						10'd619	:	dt	<=	106	;
						10'd620	:	dt	<=	101	;
						10'd621	:	dt	<=	95	;
						10'd622	:	dt	<=	86	;
						10'd623	:	dt	<=	84	;
						10'd624	:	dt	<=	85	;
						10'd625	:	dt	<=	77	;
						10'd626	:	dt	<=	78	;
						10'd627	:	dt	<=	74	;
						10'd628	:	dt	<=	76	;
						10'd629	:	dt	<=	103	;
						10'd630	:	dt	<=	152	;
						10'd631	:	dt	<=	179	;
						10'd632	:	dt	<=	170	;
						10'd633	:	dt	<=	157	;
						10'd634	:	dt	<=	155	;
						10'd635	:	dt	<=	151	;
						10'd636	:	dt	<=	140	;
						10'd637	:	dt	<=	129	;
						10'd638	:	dt	<=	126	;
						10'd639	:	dt	<=	126	;
						10'd640	:	dt	<=	133	;
						10'd641	:	dt	<=	130	;
						10'd642	:	dt	<=	122	;
						10'd643	:	dt	<=	125	;
						10'd644	:	dt	<=	81	;
						10'd645	:	dt	<=	86	;
						10'd646	:	dt	<=	85	;
						10'd647	:	dt	<=	83	;
						10'd648	:	dt	<=	76	;
						10'd649	:	dt	<=	72	;
						10'd650	:	dt	<=	73	;
						10'd651	:	dt	<=	76	;
						10'd652	:	dt	<=	77	;
						10'd653	:	dt	<=	79	;
						10'd654	:	dt	<=	71	;
						10'd655	:	dt	<=	101	;
						10'd656	:	dt	<=	151	;
						10'd657	:	dt	<=	178	;
						10'd658	:	dt	<=	177	;
						10'd659	:	dt	<=	170	;
						10'd660	:	dt	<=	161	;
						10'd661	:	dt	<=	152	;
						10'd662	:	dt	<=	147	;
						10'd663	:	dt	<=	151	;
						10'd664	:	dt	<=	133	;
						10'd665	:	dt	<=	115	;
						10'd666	:	dt	<=	121	;
						10'd667	:	dt	<=	121	;
						10'd668	:	dt	<=	124	;
						10'd669	:	dt	<=	126	;
						10'd670	:	dt	<=	122	;
						10'd671	:	dt	<=	122	;
						10'd672	:	dt	<=	61	;
						10'd673	:	dt	<=	61	;
						10'd674	:	dt	<=	67	;
						10'd675	:	dt	<=	69	;
						10'd676	:	dt	<=	70	;
						10'd677	:	dt	<=	75	;
						10'd678	:	dt	<=	78	;
						10'd679	:	dt	<=	78	;
						10'd680	:	dt	<=	81	;
						10'd681	:	dt	<=	68	;
						10'd682	:	dt	<=	113	;
						10'd683	:	dt	<=	165	;
						10'd684	:	dt	<=	174	;
						10'd685	:	dt	<=	169	;
						10'd686	:	dt	<=	162	;
						10'd687	:	dt	<=	157	;
						10'd688	:	dt	<=	149	;
						10'd689	:	dt	<=	148	;
						10'd690	:	dt	<=	148	;
						10'd691	:	dt	<=	148	;
						10'd692	:	dt	<=	126	;
						10'd693	:	dt	<=	100	;
						10'd694	:	dt	<=	113	;
						10'd695	:	dt	<=	117	;
						10'd696	:	dt	<=	113	;
						10'd697	:	dt	<=	122	;
						10'd698	:	dt	<=	118	;
						10'd699	:	dt	<=	115	;
						10'd700	:	dt	<=	69	;
						10'd701	:	dt	<=	69	;
						10'd702	:	dt	<=	77	;
						10'd703	:	dt	<=	78	;
						10'd704	:	dt	<=	75	;
						10'd705	:	dt	<=	76	;
						10'd706	:	dt	<=	78	;
						10'd707	:	dt	<=	79	;
						10'd708	:	dt	<=	67	;
						10'd709	:	dt	<=	120	;
						10'd710	:	dt	<=	173	;
						10'd711	:	dt	<=	157	;
						10'd712	:	dt	<=	159	;
						10'd713	:	dt	<=	148	;
						10'd714	:	dt	<=	155	;
						10'd715	:	dt	<=	150	;
						10'd716	:	dt	<=	138	;
						10'd717	:	dt	<=	143	;
						10'd718	:	dt	<=	148	;
						10'd719	:	dt	<=	149	;
						10'd720	:	dt	<=	123	;
						10'd721	:	dt	<=	91	;
						10'd722	:	dt	<=	101	;
						10'd723	:	dt	<=	111	;
						10'd724	:	dt	<=	111	;
						10'd725	:	dt	<=	116	;
						10'd726	:	dt	<=	113	;
						10'd727	:	dt	<=	118	;
						10'd728	:	dt	<=	74	;
						10'd729	:	dt	<=	75	;
						10'd730	:	dt	<=	76	;
						10'd731	:	dt	<=	75	;
						10'd732	:	dt	<=	75	;
						10'd733	:	dt	<=	76	;
						10'd734	:	dt	<=	75	;
						10'd735	:	dt	<=	68	;
						10'd736	:	dt	<=	124	;
						10'd737	:	dt	<=	172	;
						10'd738	:	dt	<=	152	;
						10'd739	:	dt	<=	146	;
						10'd740	:	dt	<=	146	;
						10'd741	:	dt	<=	146	;
						10'd742	:	dt	<=	152	;
						10'd743	:	dt	<=	142	;
						10'd744	:	dt	<=	131	;
						10'd745	:	dt	<=	134	;
						10'd746	:	dt	<=	144	;
						10'd747	:	dt	<=	147	;
						10'd748	:	dt	<=	125	;
						10'd749	:	dt	<=	87	;
						10'd750	:	dt	<=	87	;
						10'd751	:	dt	<=	103	;
						10'd752	:	dt	<=	107	;
						10'd753	:	dt	<=	110	;
						10'd754	:	dt	<=	116	;
						10'd755	:	dt	<=	113	;
						10'd756	:	dt	<=	75	;
						10'd757	:	dt	<=	74	;
						10'd758	:	dt	<=	74	;
						10'd759	:	dt	<=	74	;
						10'd760	:	dt	<=	76	;
						10'd761	:	dt	<=	74	;
						10'd762	:	dt	<=	82	;
						10'd763	:	dt	<=	134	;
						10'd764	:	dt	<=	168	;
						10'd765	:	dt	<=	155	;
						10'd766	:	dt	<=	146	;
						10'd767	:	dt	<=	137	;
						10'd768	:	dt	<=	145	;
						10'd769	:	dt	<=	146	;
						10'd770	:	dt	<=	149	;
						10'd771	:	dt	<=	135	;
						10'd772	:	dt	<=	124	;
						10'd773	:	dt	<=	125	;
						10'd774	:	dt	<=	138	;
						10'd775	:	dt	<=	148	;
						10'd776	:	dt	<=	127	;
						10'd777	:	dt	<=	89	;
						10'd778	:	dt	<=	82	;
						10'd779	:	dt	<=	96	;
						10'd780	:	dt	<=	106	;
						10'd781	:	dt	<=	112	;
						10'd782	:	dt	<=	120	;
						10'd783	:	dt	<=	107	;
					endcase
				end
				5'd7	:	begin
					case (cnt)			
						10'd0	:	dt	<=	171	;
						10'd1	:	dt	<=	172	;
						10'd2	:	dt	<=	172	;
						10'd3	:	dt	<=	173	;
						10'd4	:	dt	<=	173	;
						10'd5	:	dt	<=	173	;
						10'd6	:	dt	<=	173	;
						10'd7	:	dt	<=	173	;
						10'd8	:	dt	<=	172	;
						10'd9	:	dt	<=	172	;
						10'd10	:	dt	<=	172	;
						10'd11	:	dt	<=	171	;
						10'd12	:	dt	<=	170	;
						10'd13	:	dt	<=	170	;
						10'd14	:	dt	<=	169	;
						10'd15	:	dt	<=	168	;
						10'd16	:	dt	<=	168	;
						10'd17	:	dt	<=	166	;
						10'd18	:	dt	<=	165	;
						10'd19	:	dt	<=	165	;
						10'd20	:	dt	<=	164	;
						10'd21	:	dt	<=	164	;
						10'd22	:	dt	<=	152	;
						10'd23	:	dt	<=	86	;
						10'd24	:	dt	<=	72	;
						10'd25	:	dt	<=	61	;
						10'd26	:	dt	<=	65	;
						10'd27	:	dt	<=	85	;
						10'd28	:	dt	<=	174	;
						10'd29	:	dt	<=	174	;
						10'd30	:	dt	<=	174	;
						10'd31	:	dt	<=	175	;
						10'd32	:	dt	<=	175	;
						10'd33	:	dt	<=	175	;
						10'd34	:	dt	<=	175	;
						10'd35	:	dt	<=	175	;
						10'd36	:	dt	<=	175	;
						10'd37	:	dt	<=	174	;
						10'd38	:	dt	<=	174	;
						10'd39	:	dt	<=	173	;
						10'd40	:	dt	<=	172	;
						10'd41	:	dt	<=	172	;
						10'd42	:	dt	<=	172	;
						10'd43	:	dt	<=	171	;
						10'd44	:	dt	<=	170	;
						10'd45	:	dt	<=	167	;
						10'd46	:	dt	<=	166	;
						10'd47	:	dt	<=	166	;
						10'd48	:	dt	<=	166	;
						10'd49	:	dt	<=	165	;
						10'd50	:	dt	<=	168	;
						10'd51	:	dt	<=	104	;
						10'd52	:	dt	<=	64	;
						10'd53	:	dt	<=	49	;
						10'd54	:	dt	<=	59	;
						10'd55	:	dt	<=	73	;
						10'd56	:	dt	<=	175	;
						10'd57	:	dt	<=	176	;
						10'd58	:	dt	<=	176	;
						10'd59	:	dt	<=	178	;
						10'd60	:	dt	<=	179	;
						10'd61	:	dt	<=	178	;
						10'd62	:	dt	<=	176	;
						10'd63	:	dt	<=	177	;
						10'd64	:	dt	<=	177	;
						10'd65	:	dt	<=	177	;
						10'd66	:	dt	<=	176	;
						10'd67	:	dt	<=	175	;
						10'd68	:	dt	<=	174	;
						10'd69	:	dt	<=	174	;
						10'd70	:	dt	<=	173	;
						10'd71	:	dt	<=	172	;
						10'd72	:	dt	<=	172	;
						10'd73	:	dt	<=	170	;
						10'd74	:	dt	<=	169	;
						10'd75	:	dt	<=	169	;
						10'd76	:	dt	<=	168	;
						10'd77	:	dt	<=	168	;
						10'd78	:	dt	<=	171	;
						10'd79	:	dt	<=	129	;
						10'd80	:	dt	<=	49	;
						10'd81	:	dt	<=	38	;
						10'd82	:	dt	<=	56	;
						10'd83	:	dt	<=	63	;
						10'd84	:	dt	<=	178	;
						10'd85	:	dt	<=	179	;
						10'd86	:	dt	<=	181	;
						10'd87	:	dt	<=	180	;
						10'd88	:	dt	<=	181	;
						10'd89	:	dt	<=	181	;
						10'd90	:	dt	<=	180	;
						10'd91	:	dt	<=	179	;
						10'd92	:	dt	<=	179	;
						10'd93	:	dt	<=	179	;
						10'd94	:	dt	<=	178	;
						10'd95	:	dt	<=	178	;
						10'd96	:	dt	<=	178	;
						10'd97	:	dt	<=	177	;
						10'd98	:	dt	<=	175	;
						10'd99	:	dt	<=	174	;
						10'd100	:	dt	<=	174	;
						10'd101	:	dt	<=	173	;
						10'd102	:	dt	<=	172	;
						10'd103	:	dt	<=	171	;
						10'd104	:	dt	<=	170	;
						10'd105	:	dt	<=	169	;
						10'd106	:	dt	<=	169	;
						10'd107	:	dt	<=	159	;
						10'd108	:	dt	<=	59	;
						10'd109	:	dt	<=	32	;
						10'd110	:	dt	<=	44	;
						10'd111	:	dt	<=	57	;
						10'd112	:	dt	<=	179	;
						10'd113	:	dt	<=	180	;
						10'd114	:	dt	<=	182	;
						10'd115	:	dt	<=	181	;
						10'd116	:	dt	<=	182	;
						10'd117	:	dt	<=	181	;
						10'd118	:	dt	<=	181	;
						10'd119	:	dt	<=	181	;
						10'd120	:	dt	<=	181	;
						10'd121	:	dt	<=	181	;
						10'd122	:	dt	<=	180	;
						10'd123	:	dt	<=	180	;
						10'd124	:	dt	<=	180	;
						10'd125	:	dt	<=	180	;
						10'd126	:	dt	<=	177	;
						10'd127	:	dt	<=	176	;
						10'd128	:	dt	<=	176	;
						10'd129	:	dt	<=	175	;
						10'd130	:	dt	<=	173	;
						10'd131	:	dt	<=	172	;
						10'd132	:	dt	<=	172	;
						10'd133	:	dt	<=	170	;
						10'd134	:	dt	<=	170	;
						10'd135	:	dt	<=	171	;
						10'd136	:	dt	<=	122	;
						10'd137	:	dt	<=	71	;
						10'd138	:	dt	<=	53	;
						10'd139	:	dt	<=	71	;
						10'd140	:	dt	<=	180	;
						10'd141	:	dt	<=	181	;
						10'd142	:	dt	<=	182	;
						10'd143	:	dt	<=	183	;
						10'd144	:	dt	<=	184	;
						10'd145	:	dt	<=	182	;
						10'd146	:	dt	<=	183	;
						10'd147	:	dt	<=	184	;
						10'd148	:	dt	<=	184	;
						10'd149	:	dt	<=	183	;
						10'd150	:	dt	<=	181	;
						10'd151	:	dt	<=	181	;
						10'd152	:	dt	<=	180	;
						10'd153	:	dt	<=	169	;
						10'd154	:	dt	<=	168	;
						10'd155	:	dt	<=	172	;
						10'd156	:	dt	<=	171	;
						10'd157	:	dt	<=	164	;
						10'd158	:	dt	<=	158	;
						10'd159	:	dt	<=	161	;
						10'd160	:	dt	<=	153	;
						10'd161	:	dt	<=	169	;
						10'd162	:	dt	<=	168	;
						10'd163	:	dt	<=	166	;
						10'd164	:	dt	<=	128	;
						10'd165	:	dt	<=	132	;
						10'd166	:	dt	<=	142	;
						10'd167	:	dt	<=	130	;
						10'd168	:	dt	<=	182	;
						10'd169	:	dt	<=	184	;
						10'd170	:	dt	<=	185	;
						10'd171	:	dt	<=	186	;
						10'd172	:	dt	<=	187	;
						10'd173	:	dt	<=	186	;
						10'd174	:	dt	<=	186	;
						10'd175	:	dt	<=	185	;
						10'd176	:	dt	<=	184	;
						10'd177	:	dt	<=	184	;
						10'd178	:	dt	<=	183	;
						10'd179	:	dt	<=	185	;
						10'd180	:	dt	<=	183	;
						10'd181	:	dt	<=	163	;
						10'd182	:	dt	<=	152	;
						10'd183	:	dt	<=	171	;
						10'd184	:	dt	<=	176	;
						10'd185	:	dt	<=	163	;
						10'd186	:	dt	<=	151	;
						10'd187	:	dt	<=	151	;
						10'd188	:	dt	<=	140	;
						10'd189	:	dt	<=	175	;
						10'd190	:	dt	<=	164	;
						10'd191	:	dt	<=	151	;
						10'd192	:	dt	<=	94	;
						10'd193	:	dt	<=	155	;
						10'd194	:	dt	<=	166	;
						10'd195	:	dt	<=	158	;
						10'd196	:	dt	<=	185	;
						10'd197	:	dt	<=	187	;
						10'd198	:	dt	<=	188	;
						10'd199	:	dt	<=	188	;
						10'd200	:	dt	<=	187	;
						10'd201	:	dt	<=	187	;
						10'd202	:	dt	<=	188	;
						10'd203	:	dt	<=	188	;
						10'd204	:	dt	<=	189	;
						10'd205	:	dt	<=	195	;
						10'd206	:	dt	<=	200	;
						10'd207	:	dt	<=	198	;
						10'd208	:	dt	<=	187	;
						10'd209	:	dt	<=	166	;
						10'd210	:	dt	<=	159	;
						10'd211	:	dt	<=	165	;
						10'd212	:	dt	<=	152	;
						10'd213	:	dt	<=	151	;
						10'd214	:	dt	<=	136	;
						10'd215	:	dt	<=	134	;
						10'd216	:	dt	<=	129	;
						10'd217	:	dt	<=	127	;
						10'd218	:	dt	<=	128	;
						10'd219	:	dt	<=	156	;
						10'd220	:	dt	<=	114	;
						10'd221	:	dt	<=	163	;
						10'd222	:	dt	<=	127	;
						10'd223	:	dt	<=	148	;
						10'd224	:	dt	<=	186	;
						10'd225	:	dt	<=	188	;
						10'd226	:	dt	<=	188	;
						10'd227	:	dt	<=	190	;
						10'd228	:	dt	<=	189	;
						10'd229	:	dt	<=	186	;
						10'd230	:	dt	<=	184	;
						10'd231	:	dt	<=	193	;
						10'd232	:	dt	<=	203	;
						10'd233	:	dt	<=	206	;
						10'd234	:	dt	<=	205	;
						10'd235	:	dt	<=	195	;
						10'd236	:	dt	<=	185	;
						10'd237	:	dt	<=	176	;
						10'd238	:	dt	<=	175	;
						10'd239	:	dt	<=	165	;
						10'd240	:	dt	<=	129	;
						10'd241	:	dt	<=	128	;
						10'd242	:	dt	<=	152	;
						10'd243	:	dt	<=	141	;
						10'd244	:	dt	<=	135	;
						10'd245	:	dt	<=	125	;
						10'd246	:	dt	<=	122	;
						10'd247	:	dt	<=	124	;
						10'd248	:	dt	<=	112	;
						10'd249	:	dt	<=	138	;
						10'd250	:	dt	<=	114	;
						10'd251	:	dt	<=	172	;
						10'd252	:	dt	<=	187	;
						10'd253	:	dt	<=	190	;
						10'd254	:	dt	<=	191	;
						10'd255	:	dt	<=	191	;
						10'd256	:	dt	<=	206	;
						10'd257	:	dt	<=	197	;
						10'd258	:	dt	<=	187	;
						10'd259	:	dt	<=	189	;
						10'd260	:	dt	<=	196	;
						10'd261	:	dt	<=	195	;
						10'd262	:	dt	<=	191	;
						10'd263	:	dt	<=	188	;
						10'd264	:	dt	<=	186	;
						10'd265	:	dt	<=	185	;
						10'd266	:	dt	<=	179	;
						10'd267	:	dt	<=	161	;
						10'd268	:	dt	<=	142	;
						10'd269	:	dt	<=	134	;
						10'd270	:	dt	<=	150	;
						10'd271	:	dt	<=	147	;
						10'd272	:	dt	<=	140	;
						10'd273	:	dt	<=	139	;
						10'd274	:	dt	<=	124	;
						10'd275	:	dt	<=	105	;
						10'd276	:	dt	<=	106	;
						10'd277	:	dt	<=	138	;
						10'd278	:	dt	<=	122	;
						10'd279	:	dt	<=	176	;
						10'd280	:	dt	<=	189	;
						10'd281	:	dt	<=	191	;
						10'd282	:	dt	<=	190	;
						10'd283	:	dt	<=	204	;
						10'd284	:	dt	<=	220	;
						10'd285	:	dt	<=	206	;
						10'd286	:	dt	<=	193	;
						10'd287	:	dt	<=	186	;
						10'd288	:	dt	<=	190	;
						10'd289	:	dt	<=	193	;
						10'd290	:	dt	<=	191	;
						10'd291	:	dt	<=	190	;
						10'd292	:	dt	<=	188	;
						10'd293	:	dt	<=	183	;
						10'd294	:	dt	<=	179	;
						10'd295	:	dt	<=	156	;
						10'd296	:	dt	<=	143	;
						10'd297	:	dt	<=	135	;
						10'd298	:	dt	<=	126	;
						10'd299	:	dt	<=	118	;
						10'd300	:	dt	<=	115	;
						10'd301	:	dt	<=	114	;
						10'd302	:	dt	<=	103	;
						10'd303	:	dt	<=	96	;
						10'd304	:	dt	<=	89	;
						10'd305	:	dt	<=	102	;
						10'd306	:	dt	<=	126	;
						10'd307	:	dt	<=	164	;
						10'd308	:	dt	<=	190	;
						10'd309	:	dt	<=	191	;
						10'd310	:	dt	<=	192	;
						10'd311	:	dt	<=	220	;
						10'd312	:	dt	<=	221	;
						10'd313	:	dt	<=	206	;
						10'd314	:	dt	<=	178	;
						10'd315	:	dt	<=	169	;
						10'd316	:	dt	<=	179	;
						10'd317	:	dt	<=	190	;
						10'd318	:	dt	<=	190	;
						10'd319	:	dt	<=	186	;
						10'd320	:	dt	<=	178	;
						10'd321	:	dt	<=	165	;
						10'd322	:	dt	<=	153	;
						10'd323	:	dt	<=	133	;
						10'd324	:	dt	<=	120	;
						10'd325	:	dt	<=	112	;
						10'd326	:	dt	<=	108	;
						10'd327	:	dt	<=	112	;
						10'd328	:	dt	<=	117	;
						10'd329	:	dt	<=	125	;
						10'd330	:	dt	<=	123	;
						10'd331	:	dt	<=	130	;
						10'd332	:	dt	<=	140	;
						10'd333	:	dt	<=	150	;
						10'd334	:	dt	<=	169	;
						10'd335	:	dt	<=	175	;
						10'd336	:	dt	<=	193	;
						10'd337	:	dt	<=	193	;
						10'd338	:	dt	<=	202	;
						10'd339	:	dt	<=	226	;
						10'd340	:	dt	<=	217	;
						10'd341	:	dt	<=	197	;
						10'd342	:	dt	<=	166	;
						10'd343	:	dt	<=	167	;
						10'd344	:	dt	<=	177	;
						10'd345	:	dt	<=	169	;
						10'd346	:	dt	<=	163	;
						10'd347	:	dt	<=	153	;
						10'd348	:	dt	<=	141	;
						10'd349	:	dt	<=	132	;
						10'd350	:	dt	<=	120	;
						10'd351	:	dt	<=	106	;
						10'd352	:	dt	<=	105	;
						10'd353	:	dt	<=	163	;
						10'd354	:	dt	<=	184	;
						10'd355	:	dt	<=	181	;
						10'd356	:	dt	<=	183	;
						10'd357	:	dt	<=	184	;
						10'd358	:	dt	<=	182	;
						10'd359	:	dt	<=	183	;
						10'd360	:	dt	<=	181	;
						10'd361	:	dt	<=	180	;
						10'd362	:	dt	<=	168	;
						10'd363	:	dt	<=	116	;
						10'd364	:	dt	<=	195	;
						10'd365	:	dt	<=	193	;
						10'd366	:	dt	<=	218	;
						10'd367	:	dt	<=	224	;
						10'd368	:	dt	<=	213	;
						10'd369	:	dt	<=	193	;
						10'd370	:	dt	<=	182	;
						10'd371	:	dt	<=	176	;
						10'd372	:	dt	<=	163	;
						10'd373	:	dt	<=	154	;
						10'd374	:	dt	<=	158	;
						10'd375	:	dt	<=	162	;
						10'd376	:	dt	<=	156	;
						10'd377	:	dt	<=	150	;
						10'd378	:	dt	<=	145	;
						10'd379	:	dt	<=	148	;
						10'd380	:	dt	<=	129	;
						10'd381	:	dt	<=	99	;
						10'd382	:	dt	<=	166	;
						10'd383	:	dt	<=	191	;
						10'd384	:	dt	<=	188	;
						10'd385	:	dt	<=	185	;
						10'd386	:	dt	<=	184	;
						10'd387	:	dt	<=	182	;
						10'd388	:	dt	<=	180	;
						10'd389	:	dt	<=	179	;
						10'd390	:	dt	<=	178	;
						10'd391	:	dt	<=	121	;
						10'd392	:	dt	<=	193	;
						10'd393	:	dt	<=	201	;
						10'd394	:	dt	<=	229	;
						10'd395	:	dt	<=	222	;
						10'd396	:	dt	<=	218	;
						10'd397	:	dt	<=	215	;
						10'd398	:	dt	<=	211	;
						10'd399	:	dt	<=	185	;
						10'd400	:	dt	<=	162	;
						10'd401	:	dt	<=	166	;
						10'd402	:	dt	<=	167	;
						10'd403	:	dt	<=	166	;
						10'd404	:	dt	<=	156	;
						10'd405	:	dt	<=	146	;
						10'd406	:	dt	<=	142	;
						10'd407	:	dt	<=	139	;
						10'd408	:	dt	<=	120	;
						10'd409	:	dt	<=	67	;
						10'd410	:	dt	<=	58	;
						10'd411	:	dt	<=	174	;
						10'd412	:	dt	<=	190	;
						10'd413	:	dt	<=	186	;
						10'd414	:	dt	<=	184	;
						10'd415	:	dt	<=	184	;
						10'd416	:	dt	<=	181	;
						10'd417	:	dt	<=	180	;
						10'd418	:	dt	<=	179	;
						10'd419	:	dt	<=	164	;
						10'd420	:	dt	<=	190	;
						10'd421	:	dt	<=	217	;
						10'd422	:	dt	<=	228	;
						10'd423	:	dt	<=	225	;
						10'd424	:	dt	<=	223	;
						10'd425	:	dt	<=	223	;
						10'd426	:	dt	<=	218	;
						10'd427	:	dt	<=	180	;
						10'd428	:	dt	<=	148	;
						10'd429	:	dt	<=	158	;
						10'd430	:	dt	<=	156	;
						10'd431	:	dt	<=	150	;
						10'd432	:	dt	<=	143	;
						10'd433	:	dt	<=	139	;
						10'd434	:	dt	<=	132	;
						10'd435	:	dt	<=	122	;
						10'd436	:	dt	<=	105	;
						10'd437	:	dt	<=	72	;
						10'd438	:	dt	<=	41	;
						10'd439	:	dt	<=	150	;
						10'd440	:	dt	<=	193	;
						10'd441	:	dt	<=	188	;
						10'd442	:	dt	<=	186	;
						10'd443	:	dt	<=	184	;
						10'd444	:	dt	<=	183	;
						10'd445	:	dt	<=	180	;
						10'd446	:	dt	<=	179	;
						10'd447	:	dt	<=	179	;
						10'd448	:	dt	<=	205	;
						10'd449	:	dt	<=	229	;
						10'd450	:	dt	<=	228	;
						10'd451	:	dt	<=	225	;
						10'd452	:	dt	<=	222	;
						10'd453	:	dt	<=	218	;
						10'd454	:	dt	<=	206	;
						10'd455	:	dt	<=	172	;
						10'd456	:	dt	<=	152	;
						10'd457	:	dt	<=	139	;
						10'd458	:	dt	<=	117	;
						10'd459	:	dt	<=	104	;
						10'd460	:	dt	<=	113	;
						10'd461	:	dt	<=	127	;
						10'd462	:	dt	<=	137	;
						10'd463	:	dt	<=	143	;
						10'd464	:	dt	<=	143	;
						10'd465	:	dt	<=	85	;
						10'd466	:	dt	<=	69	;
						10'd467	:	dt	<=	175	;
						10'd468	:	dt	<=	191	;
						10'd469	:	dt	<=	188	;
						10'd470	:	dt	<=	188	;
						10'd471	:	dt	<=	186	;
						10'd472	:	dt	<=	185	;
						10'd473	:	dt	<=	182	;
						10'd474	:	dt	<=	181	;
						10'd475	:	dt	<=	178	;
						10'd476	:	dt	<=	226	;
						10'd477	:	dt	<=	230	;
						10'd478	:	dt	<=	229	;
						10'd479	:	dt	<=	226	;
						10'd480	:	dt	<=	220	;
						10'd481	:	dt	<=	211	;
						10'd482	:	dt	<=	197	;
						10'd483	:	dt	<=	178	;
						10'd484	:	dt	<=	160	;
						10'd485	:	dt	<=	143	;
						10'd486	:	dt	<=	123	;
						10'd487	:	dt	<=	124	;
						10'd488	:	dt	<=	154	;
						10'd489	:	dt	<=	170	;
						10'd490	:	dt	<=	158	;
						10'd491	:	dt	<=	147	;
						10'd492	:	dt	<=	156	;
						10'd493	:	dt	<=	108	;
						10'd494	:	dt	<=	169	;
						10'd495	:	dt	<=	193	;
						10'd496	:	dt	<=	190	;
						10'd497	:	dt	<=	189	;
						10'd498	:	dt	<=	189	;
						10'd499	:	dt	<=	187	;
						10'd500	:	dt	<=	185	;
						10'd501	:	dt	<=	184	;
						10'd502	:	dt	<=	181	;
						10'd503	:	dt	<=	179	;
						10'd504	:	dt	<=	228	;
						10'd505	:	dt	<=	230	;
						10'd506	:	dt	<=	229	;
						10'd507	:	dt	<=	224	;
						10'd508	:	dt	<=	214	;
						10'd509	:	dt	<=	205	;
						10'd510	:	dt	<=	188	;
						10'd511	:	dt	<=	167	;
						10'd512	:	dt	<=	165	;
						10'd513	:	dt	<=	165	;
						10'd514	:	dt	<=	145	;
						10'd515	:	dt	<=	152	;
						10'd516	:	dt	<=	164	;
						10'd517	:	dt	<=	155	;
						10'd518	:	dt	<=	145	;
						10'd519	:	dt	<=	135	;
						10'd520	:	dt	<=	129	;
						10'd521	:	dt	<=	96	;
						10'd522	:	dt	<=	186	;
						10'd523	:	dt	<=	195	;
						10'd524	:	dt	<=	192	;
						10'd525	:	dt	<=	191	;
						10'd526	:	dt	<=	190	;
						10'd527	:	dt	<=	188	;
						10'd528	:	dt	<=	186	;
						10'd529	:	dt	<=	184	;
						10'd530	:	dt	<=	183	;
						10'd531	:	dt	<=	181	;
						10'd532	:	dt	<=	229	;
						10'd533	:	dt	<=	229	;
						10'd534	:	dt	<=	226	;
						10'd535	:	dt	<=	221	;
						10'd536	:	dt	<=	208	;
						10'd537	:	dt	<=	187	;
						10'd538	:	dt	<=	165	;
						10'd539	:	dt	<=	172	;
						10'd540	:	dt	<=	187	;
						10'd541	:	dt	<=	176	;
						10'd542	:	dt	<=	154	;
						10'd543	:	dt	<=	152	;
						10'd544	:	dt	<=	148	;
						10'd545	:	dt	<=	138	;
						10'd546	:	dt	<=	132	;
						10'd547	:	dt	<=	122	;
						10'd548	:	dt	<=	101	;
						10'd549	:	dt	<=	91	;
						10'd550	:	dt	<=	192	;
						10'd551	:	dt	<=	196	;
						10'd552	:	dt	<=	194	;
						10'd553	:	dt	<=	192	;
						10'd554	:	dt	<=	190	;
						10'd555	:	dt	<=	190	;
						10'd556	:	dt	<=	188	;
						10'd557	:	dt	<=	186	;
						10'd558	:	dt	<=	184	;
						10'd559	:	dt	<=	182	;
						10'd560	:	dt	<=	230	;
						10'd561	:	dt	<=	227	;
						10'd562	:	dt	<=	223	;
						10'd563	:	dt	<=	215	;
						10'd564	:	dt	<=	196	;
						10'd565	:	dt	<=	183	;
						10'd566	:	dt	<=	185	;
						10'd567	:	dt	<=	199	;
						10'd568	:	dt	<=	197	;
						10'd569	:	dt	<=	180	;
						10'd570	:	dt	<=	157	;
						10'd571	:	dt	<=	130	;
						10'd572	:	dt	<=	117	;
						10'd573	:	dt	<=	105	;
						10'd574	:	dt	<=	92	;
						10'd575	:	dt	<=	80	;
						10'd576	:	dt	<=	83	;
						10'd577	:	dt	<=	153	;
						10'd578	:	dt	<=	199	;
						10'd579	:	dt	<=	196	;
						10'd580	:	dt	<=	196	;
						10'd581	:	dt	<=	194	;
						10'd582	:	dt	<=	192	;
						10'd583	:	dt	<=	190	;
						10'd584	:	dt	<=	189	;
						10'd585	:	dt	<=	188	;
						10'd586	:	dt	<=	185	;
						10'd587	:	dt	<=	182	;
						10'd588	:	dt	<=	227	;
						10'd589	:	dt	<=	221	;
						10'd590	:	dt	<=	214	;
						10'd591	:	dt	<=	204	;
						10'd592	:	dt	<=	197	;
						10'd593	:	dt	<=	197	;
						10'd594	:	dt	<=	199	;
						10'd595	:	dt	<=	195	;
						10'd596	:	dt	<=	186	;
						10'd597	:	dt	<=	163	;
						10'd598	:	dt	<=	132	;
						10'd599	:	dt	<=	105	;
						10'd600	:	dt	<=	101	;
						10'd601	:	dt	<=	114	;
						10'd602	:	dt	<=	90	;
						10'd603	:	dt	<=	131	;
						10'd604	:	dt	<=	178	;
						10'd605	:	dt	<=	199	;
						10'd606	:	dt	<=	198	;
						10'd607	:	dt	<=	197	;
						10'd608	:	dt	<=	196	;
						10'd609	:	dt	<=	195	;
						10'd610	:	dt	<=	193	;
						10'd611	:	dt	<=	190	;
						10'd612	:	dt	<=	188	;
						10'd613	:	dt	<=	188	;
						10'd614	:	dt	<=	185	;
						10'd615	:	dt	<=	184	;
						10'd616	:	dt	<=	219	;
						10'd617	:	dt	<=	212	;
						10'd618	:	dt	<=	206	;
						10'd619	:	dt	<=	203	;
						10'd620	:	dt	<=	203	;
						10'd621	:	dt	<=	202	;
						10'd622	:	dt	<=	188	;
						10'd623	:	dt	<=	178	;
						10'd624	:	dt	<=	173	;
						10'd625	:	dt	<=	152	;
						10'd626	:	dt	<=	124	;
						10'd627	:	dt	<=	107	;
						10'd628	:	dt	<=	173	;
						10'd629	:	dt	<=	203	;
						10'd630	:	dt	<=	196	;
						10'd631	:	dt	<=	203	;
						10'd632	:	dt	<=	203	;
						10'd633	:	dt	<=	200	;
						10'd634	:	dt	<=	200	;
						10'd635	:	dt	<=	197	;
						10'd636	:	dt	<=	196	;
						10'd637	:	dt	<=	196	;
						10'd638	:	dt	<=	194	;
						10'd639	:	dt	<=	193	;
						10'd640	:	dt	<=	189	;
						10'd641	:	dt	<=	188	;
						10'd642	:	dt	<=	187	;
						10'd643	:	dt	<=	186	;
						10'd644	:	dt	<=	207	;
						10'd645	:	dt	<=	205	;
						10'd646	:	dt	<=	207	;
						10'd647	:	dt	<=	200	;
						10'd648	:	dt	<=	196	;
						10'd649	:	dt	<=	194	;
						10'd650	:	dt	<=	180	;
						10'd651	:	dt	<=	175	;
						10'd652	:	dt	<=	162	;
						10'd653	:	dt	<=	128	;
						10'd654	:	dt	<=	100	;
						10'd655	:	dt	<=	175	;
						10'd656	:	dt	<=	209	;
						10'd657	:	dt	<=	205	;
						10'd658	:	dt	<=	205	;
						10'd659	:	dt	<=	203	;
						10'd660	:	dt	<=	201	;
						10'd661	:	dt	<=	201	;
						10'd662	:	dt	<=	200	;
						10'd663	:	dt	<=	199	;
						10'd664	:	dt	<=	197	;
						10'd665	:	dt	<=	196	;
						10'd666	:	dt	<=	195	;
						10'd667	:	dt	<=	194	;
						10'd668	:	dt	<=	192	;
						10'd669	:	dt	<=	190	;
						10'd670	:	dt	<=	188	;
						10'd671	:	dt	<=	185	;
						10'd672	:	dt	<=	199	;
						10'd673	:	dt	<=	196	;
						10'd674	:	dt	<=	200	;
						10'd675	:	dt	<=	194	;
						10'd676	:	dt	<=	185	;
						10'd677	:	dt	<=	181	;
						10'd678	:	dt	<=	174	;
						10'd679	:	dt	<=	158	;
						10'd680	:	dt	<=	126	;
						10'd681	:	dt	<=	95	;
						10'd682	:	dt	<=	164	;
						10'd683	:	dt	<=	210	;
						10'd684	:	dt	<=	206	;
						10'd685	:	dt	<=	205	;
						10'd686	:	dt	<=	203	;
						10'd687	:	dt	<=	202	;
						10'd688	:	dt	<=	202	;
						10'd689	:	dt	<=	202	;
						10'd690	:	dt	<=	202	;
						10'd691	:	dt	<=	199	;
						10'd692	:	dt	<=	199	;
						10'd693	:	dt	<=	197	;
						10'd694	:	dt	<=	196	;
						10'd695	:	dt	<=	194	;
						10'd696	:	dt	<=	192	;
						10'd697	:	dt	<=	190	;
						10'd698	:	dt	<=	189	;
						10'd699	:	dt	<=	180	;
						10'd700	:	dt	<=	198	;
						10'd701	:	dt	<=	192	;
						10'd702	:	dt	<=	187	;
						10'd703	:	dt	<=	177	;
						10'd704	:	dt	<=	167	;
						10'd705	:	dt	<=	164	;
						10'd706	:	dt	<=	151	;
						10'd707	:	dt	<=	124	;
						10'd708	:	dt	<=	92	;
						10'd709	:	dt	<=	152	;
						10'd710	:	dt	<=	210	;
						10'd711	:	dt	<=	206	;
						10'd712	:	dt	<=	204	;
						10'd713	:	dt	<=	204	;
						10'd714	:	dt	<=	203	;
						10'd715	:	dt	<=	202	;
						10'd716	:	dt	<=	201	;
						10'd717	:	dt	<=	201	;
						10'd718	:	dt	<=	199	;
						10'd719	:	dt	<=	197	;
						10'd720	:	dt	<=	197	;
						10'd721	:	dt	<=	196	;
						10'd722	:	dt	<=	196	;
						10'd723	:	dt	<=	194	;
						10'd724	:	dt	<=	192	;
						10'd725	:	dt	<=	193	;
						10'd726	:	dt	<=	188	;
						10'd727	:	dt	<=	171	;
						10'd728	:	dt	<=	193	;
						10'd729	:	dt	<=	184	;
						10'd730	:	dt	<=	172	;
						10'd731	:	dt	<=	155	;
						10'd732	:	dt	<=	147	;
						10'd733	:	dt	<=	137	;
						10'd734	:	dt	<=	112	;
						10'd735	:	dt	<=	92	;
						10'd736	:	dt	<=	153	;
						10'd737	:	dt	<=	209	;
						10'd738	:	dt	<=	208	;
						10'd739	:	dt	<=	207	;
						10'd740	:	dt	<=	205	;
						10'd741	:	dt	<=	205	;
						10'd742	:	dt	<=	203	;
						10'd743	:	dt	<=	202	;
						10'd744	:	dt	<=	201	;
						10'd745	:	dt	<=	201	;
						10'd746	:	dt	<=	199	;
						10'd747	:	dt	<=	198	;
						10'd748	:	dt	<=	197	;
						10'd749	:	dt	<=	196	;
						10'd750	:	dt	<=	195	;
						10'd751	:	dt	<=	192	;
						10'd752	:	dt	<=	192	;
						10'd753	:	dt	<=	170	;
						10'd754	:	dt	<=	165	;
						10'd755	:	dt	<=	177	;
						10'd756	:	dt	<=	173	;
						10'd757	:	dt	<=	160	;
						10'd758	:	dt	<=	143	;
						10'd759	:	dt	<=	127	;
						10'd760	:	dt	<=	115	;
						10'd761	:	dt	<=	100	;
						10'd762	:	dt	<=	85	;
						10'd763	:	dt	<=	155	;
						10'd764	:	dt	<=	212	;
						10'd765	:	dt	<=	207	;
						10'd766	:	dt	<=	208	;
						10'd767	:	dt	<=	207	;
						10'd768	:	dt	<=	207	;
						10'd769	:	dt	<=	205	;
						10'd770	:	dt	<=	203	;
						10'd771	:	dt	<=	202	;
						10'd772	:	dt	<=	201	;
						10'd773	:	dt	<=	201	;
						10'd774	:	dt	<=	199	;
						10'd775	:	dt	<=	199	;
						10'd776	:	dt	<=	198	;
						10'd777	:	dt	<=	196	;
						10'd778	:	dt	<=	195	;
						10'd779	:	dt	<=	194	;
						10'd780	:	dt	<=	183	;
						10'd781	:	dt	<=	85	;
						10'd782	:	dt	<=	65	;
						10'd783	:	dt	<=	124	;		
					endcase
				end
				5'd8	:	begin
					case (cnt)
						10'd0	:	dt	<=	212	;
						10'd1	:	dt	<=	212	;
						10'd2	:	dt	<=	213	;
						10'd3	:	dt	<=	212	;
						10'd4	:	dt	<=	214	;
						10'd5	:	dt	<=	213	;
						10'd6	:	dt	<=	213	;
						10'd7	:	dt	<=	213	;
						10'd8	:	dt	<=	214	;
						10'd9	:	dt	<=	215	;
						10'd10	:	dt	<=	214	;
						10'd11	:	dt	<=	213	;
						10'd12	:	dt	<=	212	;
						10'd13	:	dt	<=	213	;
						10'd14	:	dt	<=	212	;
						10'd15	:	dt	<=	212	;
						10'd16	:	dt	<=	211	;
						10'd17	:	dt	<=	211	;
						10'd18	:	dt	<=	212	;
						10'd19	:	dt	<=	211	;
						10'd20	:	dt	<=	210	;
						10'd21	:	dt	<=	210	;
						10'd22	:	dt	<=	207	;
						10'd23	:	dt	<=	207	;
						10'd24	:	dt	<=	207	;
						10'd25	:	dt	<=	210	;
						10'd26	:	dt	<=	191	;
						10'd27	:	dt	<=	83	;
						10'd28	:	dt	<=	213	;
						10'd29	:	dt	<=	214	;
						10'd30	:	dt	<=	215	;
						10'd31	:	dt	<=	216	;
						10'd32	:	dt	<=	216	;
						10'd33	:	dt	<=	214	;
						10'd34	:	dt	<=	215	;
						10'd35	:	dt	<=	216	;
						10'd36	:	dt	<=	216	;
						10'd37	:	dt	<=	214	;
						10'd38	:	dt	<=	212	;
						10'd39	:	dt	<=	215	;
						10'd40	:	dt	<=	214	;
						10'd41	:	dt	<=	214	;
						10'd42	:	dt	<=	216	;
						10'd43	:	dt	<=	215	;
						10'd44	:	dt	<=	213	;
						10'd45	:	dt	<=	213	;
						10'd46	:	dt	<=	213	;
						10'd47	:	dt	<=	213	;
						10'd48	:	dt	<=	212	;
						10'd49	:	dt	<=	212	;
						10'd50	:	dt	<=	209	;
						10'd51	:	dt	<=	210	;
						10'd52	:	dt	<=	210	;
						10'd53	:	dt	<=	209	;
						10'd54	:	dt	<=	208	;
						10'd55	:	dt	<=	152	;
						10'd56	:	dt	<=	216	;
						10'd57	:	dt	<=	218	;
						10'd58	:	dt	<=	218	;
						10'd59	:	dt	<=	217	;
						10'd60	:	dt	<=	217	;
						10'd61	:	dt	<=	218	;
						10'd62	:	dt	<=	216	;
						10'd63	:	dt	<=	217	;
						10'd64	:	dt	<=	219	;
						10'd65	:	dt	<=	222	;
						10'd66	:	dt	<=	163	;
						10'd67	:	dt	<=	205	;
						10'd68	:	dt	<=	222	;
						10'd69	:	dt	<=	218	;
						10'd70	:	dt	<=	219	;
						10'd71	:	dt	<=	219	;
						10'd72	:	dt	<=	218	;
						10'd73	:	dt	<=	217	;
						10'd74	:	dt	<=	216	;
						10'd75	:	dt	<=	215	;
						10'd76	:	dt	<=	215	;
						10'd77	:	dt	<=	213	;
						10'd78	:	dt	<=	211	;
						10'd79	:	dt	<=	210	;
						10'd80	:	dt	<=	211	;
						10'd81	:	dt	<=	210	;
						10'd82	:	dt	<=	211	;
						10'd83	:	dt	<=	126	;
						10'd84	:	dt	<=	217	;
						10'd85	:	dt	<=	219	;
						10'd86	:	dt	<=	219	;
						10'd87	:	dt	<=	218	;
						10'd88	:	dt	<=	219	;
						10'd89	:	dt	<=	219	;
						10'd90	:	dt	<=	219	;
						10'd91	:	dt	<=	217	;
						10'd92	:	dt	<=	224	;
						10'd93	:	dt	<=	223	;
						10'd94	:	dt	<=	134	;
						10'd95	:	dt	<=	199	;
						10'd96	:	dt	<=	225	;
						10'd97	:	dt	<=	220	;
						10'd98	:	dt	<=	220	;
						10'd99	:	dt	<=	220	;
						10'd100	:	dt	<=	220	;
						10'd101	:	dt	<=	218	;
						10'd102	:	dt	<=	218	;
						10'd103	:	dt	<=	217	;
						10'd104	:	dt	<=	217	;
						10'd105	:	dt	<=	215	;
						10'd106	:	dt	<=	215	;
						10'd107	:	dt	<=	213	;
						10'd108	:	dt	<=	213	;
						10'd109	:	dt	<=	214	;
						10'd110	:	dt	<=	204	;
						10'd111	:	dt	<=	143	;
						10'd112	:	dt	<=	219	;
						10'd113	:	dt	<=	219	;
						10'd114	:	dt	<=	220	;
						10'd115	:	dt	<=	220	;
						10'd116	:	dt	<=	220	;
						10'd117	:	dt	<=	219	;
						10'd118	:	dt	<=	221	;
						10'd119	:	dt	<=	216	;
						10'd120	:	dt	<=	235	;
						10'd121	:	dt	<=	202	;
						10'd122	:	dt	<=	117	;
						10'd123	:	dt	<=	213	;
						10'd124	:	dt	<=	224	;
						10'd125	:	dt	<=	221	;
						10'd126	:	dt	<=	220	;
						10'd127	:	dt	<=	222	;
						10'd128	:	dt	<=	221	;
						10'd129	:	dt	<=	220	;
						10'd130	:	dt	<=	220	;
						10'd131	:	dt	<=	219	;
						10'd132	:	dt	<=	218	;
						10'd133	:	dt	<=	217	;
						10'd134	:	dt	<=	218	;
						10'd135	:	dt	<=	216	;
						10'd136	:	dt	<=	215	;
						10'd137	:	dt	<=	214	;
						10'd138	:	dt	<=	210	;
						10'd139	:	dt	<=	180	;
						10'd140	:	dt	<=	221	;
						10'd141	:	dt	<=	221	;
						10'd142	:	dt	<=	221	;
						10'd143	:	dt	<=	222	;
						10'd144	:	dt	<=	221	;
						10'd145	:	dt	<=	220	;
						10'd146	:	dt	<=	221	;
						10'd147	:	dt	<=	220	;
						10'd148	:	dt	<=	246	;
						10'd149	:	dt	<=	182	;
						10'd150	:	dt	<=	117	;
						10'd151	:	dt	<=	229	;
						10'd152	:	dt	<=	224	;
						10'd153	:	dt	<=	223	;
						10'd154	:	dt	<=	223	;
						10'd155	:	dt	<=	225	;
						10'd156	:	dt	<=	223	;
						10'd157	:	dt	<=	221	;
						10'd158	:	dt	<=	222	;
						10'd159	:	dt	<=	222	;
						10'd160	:	dt	<=	220	;
						10'd161	:	dt	<=	218	;
						10'd162	:	dt	<=	218	;
						10'd163	:	dt	<=	218	;
						10'd164	:	dt	<=	217	;
						10'd165	:	dt	<=	216	;
						10'd166	:	dt	<=	212	;
						10'd167	:	dt	<=	214	;
						10'd168	:	dt	<=	221	;
						10'd169	:	dt	<=	221	;
						10'd170	:	dt	<=	224	;
						10'd171	:	dt	<=	224	;
						10'd172	:	dt	<=	223	;
						10'd173	:	dt	<=	225	;
						10'd174	:	dt	<=	222	;
						10'd175	:	dt	<=	226	;
						10'd176	:	dt	<=	250	;
						10'd177	:	dt	<=	171	;
						10'd178	:	dt	<=	133	;
						10'd179	:	dt	<=	233	;
						10'd180	:	dt	<=	224	;
						10'd181	:	dt	<=	225	;
						10'd182	:	dt	<=	226	;
						10'd183	:	dt	<=	226	;
						10'd184	:	dt	<=	224	;
						10'd185	:	dt	<=	224	;
						10'd186	:	dt	<=	223	;
						10'd187	:	dt	<=	221	;
						10'd188	:	dt	<=	221	;
						10'd189	:	dt	<=	220	;
						10'd190	:	dt	<=	220	;
						10'd191	:	dt	<=	219	;
						10'd192	:	dt	<=	218	;
						10'd193	:	dt	<=	218	;
						10'd194	:	dt	<=	215	;
						10'd195	:	dt	<=	216	;
						10'd196	:	dt	<=	223	;
						10'd197	:	dt	<=	223	;
						10'd198	:	dt	<=	225	;
						10'd199	:	dt	<=	226	;
						10'd200	:	dt	<=	225	;
						10'd201	:	dt	<=	226	;
						10'd202	:	dt	<=	223	;
						10'd203	:	dt	<=	235	;
						10'd204	:	dt	<=	243	;
						10'd205	:	dt	<=	141	;
						10'd206	:	dt	<=	159	;
						10'd207	:	dt	<=	236	;
						10'd208	:	dt	<=	224	;
						10'd209	:	dt	<=	231	;
						10'd210	:	dt	<=	227	;
						10'd211	:	dt	<=	226	;
						10'd212	:	dt	<=	230	;
						10'd213	:	dt	<=	225	;
						10'd214	:	dt	<=	224	;
						10'd215	:	dt	<=	224	;
						10'd216	:	dt	<=	222	;
						10'd217	:	dt	<=	224	;
						10'd218	:	dt	<=	220	;
						10'd219	:	dt	<=	220	;
						10'd220	:	dt	<=	220	;
						10'd221	:	dt	<=	218	;
						10'd222	:	dt	<=	217	;
						10'd223	:	dt	<=	215	;
						10'd224	:	dt	<=	225	;
						10'd225	:	dt	<=	226	;
						10'd226	:	dt	<=	225	;
						10'd227	:	dt	<=	225	;
						10'd228	:	dt	<=	227	;
						10'd229	:	dt	<=	228	;
						10'd230	:	dt	<=	222	;
						10'd231	:	dt	<=	242	;
						10'd232	:	dt	<=	230	;
						10'd233	:	dt	<=	136	;
						10'd234	:	dt	<=	166	;
						10'd235	:	dt	<=	244	;
						10'd236	:	dt	<=	204	;
						10'd237	:	dt	<=	199	;
						10'd238	:	dt	<=	230	;
						10'd239	:	dt	<=	220	;
						10'd240	:	dt	<=	211	;
						10'd241	:	dt	<=	231	;
						10'd242	:	dt	<=	231	;
						10'd243	:	dt	<=	231	;
						10'd244	:	dt	<=	227	;
						10'd245	:	dt	<=	224	;
						10'd246	:	dt	<=	225	;
						10'd247	:	dt	<=	221	;
						10'd248	:	dt	<=	222	;
						10'd249	:	dt	<=	219	;
						10'd250	:	dt	<=	220	;
						10'd251	:	dt	<=	220	;
						10'd252	:	dt	<=	226	;
						10'd253	:	dt	<=	227	;
						10'd254	:	dt	<=	227	;
						10'd255	:	dt	<=	227	;
						10'd256	:	dt	<=	227	;
						10'd257	:	dt	<=	227	;
						10'd258	:	dt	<=	224	;
						10'd259	:	dt	<=	247	;
						10'd260	:	dt	<=	226	;
						10'd261	:	dt	<=	147	;
						10'd262	:	dt	<=	173	;
						10'd263	:	dt	<=	255	;
						10'd264	:	dt	<=	207	;
						10'd265	:	dt	<=	147	;
						10'd266	:	dt	<=	199	;
						10'd267	:	dt	<=	213	;
						10'd268	:	dt	<=	151	;
						10'd269	:	dt	<=	177	;
						10'd270	:	dt	<=	205	;
						10'd271	:	dt	<=	201	;
						10'd272	:	dt	<=	217	;
						10'd273	:	dt	<=	174	;
						10'd274	:	dt	<=	181	;
						10'd275	:	dt	<=	230	;
						10'd276	:	dt	<=	221	;
						10'd277	:	dt	<=	224	;
						10'd278	:	dt	<=	222	;
						10'd279	:	dt	<=	221	;
						10'd280	:	dt	<=	228	;
						10'd281	:	dt	<=	228	;
						10'd282	:	dt	<=	228	;
						10'd283	:	dt	<=	228	;
						10'd284	:	dt	<=	229	;
						10'd285	:	dt	<=	228	;
						10'd286	:	dt	<=	227	;
						10'd287	:	dt	<=	250	;
						10'd288	:	dt	<=	228	;
						10'd289	:	dt	<=	154	;
						10'd290	:	dt	<=	219	;
						10'd291	:	dt	<=	255	;
						10'd292	:	dt	<=	231	;
						10'd293	:	dt	<=	166	;
						10'd294	:	dt	<=	160	;
						10'd295	:	dt	<=	207	;
						10'd296	:	dt	<=	172	;
						10'd297	:	dt	<=	114	;
						10'd298	:	dt	<=	140	;
						10'd299	:	dt	<=	159	;
						10'd300	:	dt	<=	206	;
						10'd301	:	dt	<=	142	;
						10'd302	:	dt	<=	128	;
						10'd303	:	dt	<=	235	;
						10'd304	:	dt	<=	223	;
						10'd305	:	dt	<=	225	;
						10'd306	:	dt	<=	223	;
						10'd307	:	dt	<=	221	;
						10'd308	:	dt	<=	228	;
						10'd309	:	dt	<=	228	;
						10'd310	:	dt	<=	228	;
						10'd311	:	dt	<=	228	;
						10'd312	:	dt	<=	230	;
						10'd313	:	dt	<=	229	;
						10'd314	:	dt	<=	232	;
						10'd315	:	dt	<=	248	;
						10'd316	:	dt	<=	223	;
						10'd317	:	dt	<=	166	;
						10'd318	:	dt	<=	251	;
						10'd319	:	dt	<=	255	;
						10'd320	:	dt	<=	246	;
						10'd321	:	dt	<=	184	;
						10'd322	:	dt	<=	131	;
						10'd323	:	dt	<=	200	;
						10'd324	:	dt	<=	169	;
						10'd325	:	dt	<=	138	;
						10'd326	:	dt	<=	189	;
						10'd327	:	dt	<=	161	;
						10'd328	:	dt	<=	226	;
						10'd329	:	dt	<=	145	;
						10'd330	:	dt	<=	123	;
						10'd331	:	dt	<=	237	;
						10'd332	:	dt	<=	223	;
						10'd333	:	dt	<=	224	;
						10'd334	:	dt	<=	223	;
						10'd335	:	dt	<=	223	;
						10'd336	:	dt	<=	229	;
						10'd337	:	dt	<=	228	;
						10'd338	:	dt	<=	229	;
						10'd339	:	dt	<=	229	;
						10'd340	:	dt	<=	231	;
						10'd341	:	dt	<=	228	;
						10'd342	:	dt	<=	241	;
						10'd343	:	dt	<=	232	;
						10'd344	:	dt	<=	217	;
						10'd345	:	dt	<=	201	;
						10'd346	:	dt	<=	234	;
						10'd347	:	dt	<=	255	;
						10'd348	:	dt	<=	254	;
						10'd349	:	dt	<=	193	;
						10'd350	:	dt	<=	118	;
						10'd351	:	dt	<=	188	;
						10'd352	:	dt	<=	151	;
						10'd353	:	dt	<=	179	;
						10'd354	:	dt	<=	205	;
						10'd355	:	dt	<=	163	;
						10'd356	:	dt	<=	231	;
						10'd357	:	dt	<=	182	;
						10'd358	:	dt	<=	132	;
						10'd359	:	dt	<=	232	;
						10'd360	:	dt	<=	227	;
						10'd361	:	dt	<=	225	;
						10'd362	:	dt	<=	225	;
						10'd363	:	dt	<=	224	;
						10'd364	:	dt	<=	229	;
						10'd365	:	dt	<=	229	;
						10'd366	:	dt	<=	229	;
						10'd367	:	dt	<=	229	;
						10'd368	:	dt	<=	231	;
						10'd369	:	dt	<=	232	;
						10'd370	:	dt	<=	238	;
						10'd371	:	dt	<=	204	;
						10'd372	:	dt	<=	221	;
						10'd373	:	dt	<=	226	;
						10'd374	:	dt	<=	199	;
						10'd375	:	dt	<=	242	;
						10'd376	:	dt	<=	255	;
						10'd377	:	dt	<=	198	;
						10'd378	:	dt	<=	113	;
						10'd379	:	dt	<=	158	;
						10'd380	:	dt	<=	152	;
						10'd381	:	dt	<=	199	;
						10'd382	:	dt	<=	183	;
						10'd383	:	dt	<=	160	;
						10'd384	:	dt	<=	222	;
						10'd385	:	dt	<=	208	;
						10'd386	:	dt	<=	156	;
						10'd387	:	dt	<=	188	;
						10'd388	:	dt	<=	238	;
						10'd389	:	dt	<=	226	;
						10'd390	:	dt	<=	227	;
						10'd391	:	dt	<=	225	;
						10'd392	:	dt	<=	228	;
						10'd393	:	dt	<=	228	;
						10'd394	:	dt	<=	229	;
						10'd395	:	dt	<=	229	;
						10'd396	:	dt	<=	229	;
						10'd397	:	dt	<=	237	;
						10'd398	:	dt	<=	237	;
						10'd399	:	dt	<=	176	;
						10'd400	:	dt	<=	215	;
						10'd401	:	dt	<=	211	;
						10'd402	:	dt	<=	194	;
						10'd403	:	dt	<=	220	;
						10'd404	:	dt	<=	255	;
						10'd405	:	dt	<=	207	;
						10'd406	:	dt	<=	114	;
						10'd407	:	dt	<=	115	;
						10'd408	:	dt	<=	158	;
						10'd409	:	dt	<=	205	;
						10'd410	:	dt	<=	168	;
						10'd411	:	dt	<=	126	;
						10'd412	:	dt	<=	215	;
						10'd413	:	dt	<=	210	;
						10'd414	:	dt	<=	149	;
						10'd415	:	dt	<=	135	;
						10'd416	:	dt	<=	241	;
						10'd417	:	dt	<=	225	;
						10'd418	:	dt	<=	227	;
						10'd419	:	dt	<=	226	;
						10'd420	:	dt	<=	227	;
						10'd421	:	dt	<=	228	;
						10'd422	:	dt	<=	229	;
						10'd423	:	dt	<=	229	;
						10'd424	:	dt	<=	226	;
						10'd425	:	dt	<=	242	;
						10'd426	:	dt	<=	238	;
						10'd427	:	dt	<=	163	;
						10'd428	:	dt	<=	173	;
						10'd429	:	dt	<=	192	;
						10'd430	:	dt	<=	169	;
						10'd431	:	dt	<=	192	;
						10'd432	:	dt	<=	252	;
						10'd433	:	dt	<=	201	;
						10'd434	:	dt	<=	105	;
						10'd435	:	dt	<=	95	;
						10'd436	:	dt	<=	153	;
						10'd437	:	dt	<=	196	;
						10'd438	:	dt	<=	146	;
						10'd439	:	dt	<=	119	;
						10'd440	:	dt	<=	220	;
						10'd441	:	dt	<=	193	;
						10'd442	:	dt	<=	118	;
						10'd443	:	dt	<=	165	;
						10'd444	:	dt	<=	240	;
						10'd445	:	dt	<=	227	;
						10'd446	:	dt	<=	228	;
						10'd447	:	dt	<=	227	;
						10'd448	:	dt	<=	228	;
						10'd449	:	dt	<=	228	;
						10'd450	:	dt	<=	229	;
						10'd451	:	dt	<=	230	;
						10'd452	:	dt	<=	227	;
						10'd453	:	dt	<=	250	;
						10'd454	:	dt	<=	255	;
						10'd455	:	dt	<=	162	;
						10'd456	:	dt	<=	147	;
						10'd457	:	dt	<=	153	;
						10'd458	:	dt	<=	146	;
						10'd459	:	dt	<=	147	;
						10'd460	:	dt	<=	227	;
						10'd461	:	dt	<=	212	;
						10'd462	:	dt	<=	118	;
						10'd463	:	dt	<=	85	;
						10'd464	:	dt	<=	159	;
						10'd465	:	dt	<=	213	;
						10'd466	:	dt	<=	132	;
						10'd467	:	dt	<=	151	;
						10'd468	:	dt	<=	208	;
						10'd469	:	dt	<=	148	;
						10'd470	:	dt	<=	110	;
						10'd471	:	dt	<=	224	;
						10'd472	:	dt	<=	229	;
						10'd473	:	dt	<=	227	;
						10'd474	:	dt	<=	226	;
						10'd475	:	dt	<=	226	;
						10'd476	:	dt	<=	228	;
						10'd477	:	dt	<=	229	;
						10'd478	:	dt	<=	229	;
						10'd479	:	dt	<=	229	;
						10'd480	:	dt	<=	232	;
						10'd481	:	dt	<=	255	;
						10'd482	:	dt	<=	255	;
						10'd483	:	dt	<=	184	;
						10'd484	:	dt	<=	132	;
						10'd485	:	dt	<=	149	;
						10'd486	:	dt	<=	139	;
						10'd487	:	dt	<=	143	;
						10'd488	:	dt	<=	196	;
						10'd489	:	dt	<=	225	;
						10'd490	:	dt	<=	159	;
						10'd491	:	dt	<=	64	;
						10'd492	:	dt	<=	150	;
						10'd493	:	dt	<=	173	;
						10'd494	:	dt	<=	130	;
						10'd495	:	dt	<=	184	;
						10'd496	:	dt	<=	156	;
						10'd497	:	dt	<=	101	;
						10'd498	:	dt	<=	157	;
						10'd499	:	dt	<=	239	;
						10'd500	:	dt	<=	225	;
						10'd501	:	dt	<=	227	;
						10'd502	:	dt	<=	226	;
						10'd503	:	dt	<=	226	;
						10'd504	:	dt	<=	228	;
						10'd505	:	dt	<=	229	;
						10'd506	:	dt	<=	230	;
						10'd507	:	dt	<=	228	;
						10'd508	:	dt	<=	236	;
						10'd509	:	dt	<=	255	;
						10'd510	:	dt	<=	255	;
						10'd511	:	dt	<=	207	;
						10'd512	:	dt	<=	126	;
						10'd513	:	dt	<=	135	;
						10'd514	:	dt	<=	139	;
						10'd515	:	dt	<=	135	;
						10'd516	:	dt	<=	180	;
						10'd517	:	dt	<=	193	;
						10'd518	:	dt	<=	123	;
						10'd519	:	dt	<=	109	;
						10'd520	:	dt	<=	202	;
						10'd521	:	dt	<=	180	;
						10'd522	:	dt	<=	196	;
						10'd523	:	dt	<=	197	;
						10'd524	:	dt	<=	124	;
						10'd525	:	dt	<=	100	;
						10'd526	:	dt	<=	222	;
						10'd527	:	dt	<=	231	;
						10'd528	:	dt	<=	227	;
						10'd529	:	dt	<=	228	;
						10'd530	:	dt	<=	228	;
						10'd531	:	dt	<=	227	;
						10'd532	:	dt	<=	228	;
						10'd533	:	dt	<=	229	;
						10'd534	:	dt	<=	230	;
						10'd535	:	dt	<=	230	;
						10'd536	:	dt	<=	241	;
						10'd537	:	dt	<=	255	;
						10'd538	:	dt	<=	255	;
						10'd539	:	dt	<=	218	;
						10'd540	:	dt	<=	127	;
						10'd541	:	dt	<=	138	;
						10'd542	:	dt	<=	151	;
						10'd543	:	dt	<=	139	;
						10'd544	:	dt	<=	204	;
						10'd545	:	dt	<=	214	;
						10'd546	:	dt	<=	183	;
						10'd547	:	dt	<=	220	;
						10'd548	:	dt	<=	217	;
						10'd549	:	dt	<=	191	;
						10'd550	:	dt	<=	176	;
						10'd551	:	dt	<=	184	;
						10'd552	:	dt	<=	112	;
						10'd553	:	dt	<=	124	;
						10'd554	:	dt	<=	242	;
						10'd555	:	dt	<=	228	;
						10'd556	:	dt	<=	231	;
						10'd557	:	dt	<=	230	;
						10'd558	:	dt	<=	227	;
						10'd559	:	dt	<=	227	;
						10'd560	:	dt	<=	227	;
						10'd561	:	dt	<=	228	;
						10'd562	:	dt	<=	229	;
						10'd563	:	dt	<=	228	;
						10'd564	:	dt	<=	242	;
						10'd565	:	dt	<=	255	;
						10'd566	:	dt	<=	255	;
						10'd567	:	dt	<=	220	;
						10'd568	:	dt	<=	132	;
						10'd569	:	dt	<=	150	;
						10'd570	:	dt	<=	148	;
						10'd571	:	dt	<=	171	;
						10'd572	:	dt	<=	237	;
						10'd573	:	dt	<=	244	;
						10'd574	:	dt	<=	246	;
						10'd575	:	dt	<=	229	;
						10'd576	:	dt	<=	209	;
						10'd577	:	dt	<=	192	;
						10'd578	:	dt	<=	149	;
						10'd579	:	dt	<=	144	;
						10'd580	:	dt	<=	98	;
						10'd581	:	dt	<=	159	;
						10'd582	:	dt	<=	244	;
						10'd583	:	dt	<=	228	;
						10'd584	:	dt	<=	232	;
						10'd585	:	dt	<=	231	;
						10'd586	:	dt	<=	229	;
						10'd587	:	dt	<=	227	;
						10'd588	:	dt	<=	235	;
						10'd589	:	dt	<=	237	;
						10'd590	:	dt	<=	238	;
						10'd591	:	dt	<=	236	;
						10'd592	:	dt	<=	243	;
						10'd593	:	dt	<=	255	;
						10'd594	:	dt	<=	255	;
						10'd595	:	dt	<=	209	;
						10'd596	:	dt	<=	151	;
						10'd597	:	dt	<=	169	;
						10'd598	:	dt	<=	147	;
						10'd599	:	dt	<=	219	;
						10'd600	:	dt	<=	253	;
						10'd601	:	dt	<=	248	;
						10'd602	:	dt	<=	246	;
						10'd603	:	dt	<=	232	;
						10'd604	:	dt	<=	210	;
						10'd605	:	dt	<=	178	;
						10'd606	:	dt	<=	138	;
						10'd607	:	dt	<=	105	;
						10'd608	:	dt	<=	105	;
						10'd609	:	dt	<=	226	;
						10'd610	:	dt	<=	235	;
						10'd611	:	dt	<=	231	;
						10'd612	:	dt	<=	232	;
						10'd613	:	dt	<=	231	;
						10'd614	:	dt	<=	230	;
						10'd615	:	dt	<=	228	;
						10'd616	:	dt	<=	164	;
						10'd617	:	dt	<=	167	;
						10'd618	:	dt	<=	171	;
						10'd619	:	dt	<=	166	;
						10'd620	:	dt	<=	220	;
						10'd621	:	dt	<=	255	;
						10'd622	:	dt	<=	255	;
						10'd623	:	dt	<=	215	;
						10'd624	:	dt	<=	180	;
						10'd625	:	dt	<=	175	;
						10'd626	:	dt	<=	151	;
						10'd627	:	dt	<=	229	;
						10'd628	:	dt	<=	255	;
						10'd629	:	dt	<=	255	;
						10'd630	:	dt	<=	246	;
						10'd631	:	dt	<=	226	;
						10'd632	:	dt	<=	199	;
						10'd633	:	dt	<=	159	;
						10'd634	:	dt	<=	122	;
						10'd635	:	dt	<=	85	;
						10'd636	:	dt	<=	163	;
						10'd637	:	dt	<=	246	;
						10'd638	:	dt	<=	235	;
						10'd639	:	dt	<=	235	;
						10'd640	:	dt	<=	227	;
						10'd641	:	dt	<=	225	;
						10'd642	:	dt	<=	229	;
						10'd643	:	dt	<=	231	;
						10'd644	:	dt	<=	101	;
						10'd645	:	dt	<=	101	;
						10'd646	:	dt	<=	104	;
						10'd647	:	dt	<=	87	;
						10'd648	:	dt	<=	172	;
						10'd649	:	dt	<=	255	;
						10'd650	:	dt	<=	252	;
						10'd651	:	dt	<=	229	;
						10'd652	:	dt	<=	188	;
						10'd653	:	dt	<=	185	;
						10'd654	:	dt	<=	162	;
						10'd655	:	dt	<=	217	;
						10'd656	:	dt	<=	255	;
						10'd657	:	dt	<=	255	;
						10'd658	:	dt	<=	227	;
						10'd659	:	dt	<=	209	;
						10'd660	:	dt	<=	180	;
						10'd661	:	dt	<=	136	;
						10'd662	:	dt	<=	108	;
						10'd663	:	dt	<=	93	;
						10'd664	:	dt	<=	128	;
						10'd665	:	dt	<=	140	;
						10'd666	:	dt	<=	137	;
						10'd667	:	dt	<=	152	;
						10'd668	:	dt	<=	187	;
						10'd669	:	dt	<=	227	;
						10'd670	:	dt	<=	239	;
						10'd671	:	dt	<=	234	;
						10'd672	:	dt	<=	115	;
						10'd673	:	dt	<=	114	;
						10'd674	:	dt	<=	116	;
						10'd675	:	dt	<=	104	;
						10'd676	:	dt	<=	148	;
						10'd677	:	dt	<=	255	;
						10'd678	:	dt	<=	250	;
						10'd679	:	dt	<=	228	;
						10'd680	:	dt	<=	189	;
						10'd681	:	dt	<=	188	;
						10'd682	:	dt	<=	167	;
						10'd683	:	dt	<=	217	;
						10'd684	:	dt	<=	255	;
						10'd685	:	dt	<=	246	;
						10'd686	:	dt	<=	213	;
						10'd687	:	dt	<=	186	;
						10'd688	:	dt	<=	155	;
						10'd689	:	dt	<=	117	;
						10'd690	:	dt	<=	102	;
						10'd691	:	dt	<=	92	;
						10'd692	:	dt	<=	98	;
						10'd693	:	dt	<=	129	;
						10'd694	:	dt	<=	172	;
						10'd695	:	dt	<=	217	;
						10'd696	:	dt	<=	235	;
						10'd697	:	dt	<=	234	;
						10'd698	:	dt	<=	235	;
						10'd699	:	dt	<=	230	;
						10'd700	:	dt	<=	114	;
						10'd701	:	dt	<=	112	;
						10'd702	:	dt	<=	115	;
						10'd703	:	dt	<=	103	;
						10'd704	:	dt	<=	145	;
						10'd705	:	dt	<=	255	;
						10'd706	:	dt	<=	236	;
						10'd707	:	dt	<=	211	;
						10'd708	:	dt	<=	185	;
						10'd709	:	dt	<=	182	;
						10'd710	:	dt	<=	169	;
						10'd711	:	dt	<=	234	;
						10'd712	:	dt	<=	253	;
						10'd713	:	dt	<=	222	;
						10'd714	:	dt	<=	194	;
						10'd715	:	dt	<=	156	;
						10'd716	:	dt	<=	132	;
						10'd717	:	dt	<=	100	;
						10'd718	:	dt	<=	101	;
						10'd719	:	dt	<=	163	;
						10'd720	:	dt	<=	198	;
						10'd721	:	dt	<=	234	;
						10'd722	:	dt	<=	245	;
						10'd723	:	dt	<=	243	;
						10'd724	:	dt	<=	245	;
						10'd725	:	dt	<=	236	;
						10'd726	:	dt	<=	220	;
						10'd727	:	dt	<=	221	;
						10'd728	:	dt	<=	112	;
						10'd729	:	dt	<=	112	;
						10'd730	:	dt	<=	119	;
						10'd731	:	dt	<=	102	;
						10'd732	:	dt	<=	168	;
						10'd733	:	dt	<=	255	;
						10'd734	:	dt	<=	225	;
						10'd735	:	dt	<=	206	;
						10'd736	:	dt	<=	189	;
						10'd737	:	dt	<=	180	;
						10'd738	:	dt	<=	184	;
						10'd739	:	dt	<=	227	;
						10'd740	:	dt	<=	225	;
						10'd741	:	dt	<=	208	;
						10'd742	:	dt	<=	169	;
						10'd743	:	dt	<=	135	;
						10'd744	:	dt	<=	124	;
						10'd745	:	dt	<=	79	;
						10'd746	:	dt	<=	166	;
						10'd747	:	dt	<=	255	;
						10'd748	:	dt	<=	250	;
						10'd749	:	dt	<=	217	;
						10'd750	:	dt	<=	208	;
						10'd751	:	dt	<=	214	;
						10'd752	:	dt	<=	224	;
						10'd753	:	dt	<=	237	;
						10'd754	:	dt	<=	231	;
						10'd755	:	dt	<=	218	;
						10'd756	:	dt	<=	112	;
						10'd757	:	dt	<=	111	;
						10'd758	:	dt	<=	117	;
						10'd759	:	dt	<=	101	;
						10'd760	:	dt	<=	194	;
						10'd761	:	dt	<=	251	;
						10'd762	:	dt	<=	220	;
						10'd763	:	dt	<=	205	;
						10'd764	:	dt	<=	193	;
						10'd765	:	dt	<=	184	;
						10'd766	:	dt	<=	193	;
						10'd767	:	dt	<=	212	;
						10'd768	:	dt	<=	207	;
						10'd769	:	dt	<=	194	;
						10'd770	:	dt	<=	151	;
						10'd771	:	dt	<=	128	;
						10'd772	:	dt	<=	117	;
						10'd773	:	dt	<=	112	;
						10'd774	:	dt	<=	213	;
						10'd775	:	dt	<=	219	;
						10'd776	:	dt	<=	249	;
						10'd777	:	dt	<=	242	;
						10'd778	:	dt	<=	211	;
						10'd779	:	dt	<=	198	;
						10'd780	:	dt	<=	206	;
						10'd781	:	dt	<=	209	;
						10'd782	:	dt	<=	204	;
						10'd783	:	dt	<=	210	;
					endcase
				end
				5'd9	:	begin
				end
				5'd10	:	begin
					case (cnt)
						10'd0	:	dt	<=	93	;
						10'd1	:	dt	<=	100	;
						10'd2	:	dt	<=	112	;
						10'd3	:	dt	<=	118	;
						10'd4	:	dt	<=	123	;
						10'd5	:	dt	<=	127	;
						10'd6	:	dt	<=	131	;
						10'd7	:	dt	<=	133	;
						10'd8	:	dt	<=	136	;
						10'd9	:	dt	<=	139	;
						10'd10	:	dt	<=	140	;
						10'd11	:	dt	<=	143	;
						10'd12	:	dt	<=	144	;
						10'd13	:	dt	<=	145	;
						10'd14	:	dt	<=	146	;
						10'd15	:	dt	<=	149	;
						10'd16	:	dt	<=	151	;
						10'd17	:	dt	<=	153	;
						10'd18	:	dt	<=	154	;
						10'd19	:	dt	<=	155	;
						10'd20	:	dt	<=	156	;
						10'd21	:	dt	<=	159	;
						10'd22	:	dt	<=	159	;
						10'd23	:	dt	<=	160	;
						10'd24	:	dt	<=	160	;
						10'd25	:	dt	<=	161	;
						10'd26	:	dt	<=	163	;
						10'd27	:	dt	<=	164	;
						10'd28	:	dt	<=	93	;
						10'd29	:	dt	<=	102	;
						10'd30	:	dt	<=	113	;
						10'd31	:	dt	<=	119	;
						10'd32	:	dt	<=	123	;
						10'd33	:	dt	<=	128	;
						10'd34	:	dt	<=	131	;
						10'd35	:	dt	<=	134	;
						10'd36	:	dt	<=	138	;
						10'd37	:	dt	<=	140	;
						10'd38	:	dt	<=	141	;
						10'd39	:	dt	<=	144	;
						10'd40	:	dt	<=	145	;
						10'd41	:	dt	<=	146	;
						10'd42	:	dt	<=	148	;
						10'd43	:	dt	<=	150	;
						10'd44	:	dt	<=	137	;
						10'd45	:	dt	<=	149	;
						10'd46	:	dt	<=	155	;
						10'd47	:	dt	<=	156	;
						10'd48	:	dt	<=	158	;
						10'd49	:	dt	<=	160	;
						10'd50	:	dt	<=	160	;
						10'd51	:	dt	<=	161	;
						10'd52	:	dt	<=	162	;
						10'd53	:	dt	<=	163	;
						10'd54	:	dt	<=	164	;
						10'd55	:	dt	<=	165	;
						10'd56	:	dt	<=	95	;
						10'd57	:	dt	<=	104	;
						10'd58	:	dt	<=	114	;
						10'd59	:	dt	<=	120	;
						10'd60	:	dt	<=	124	;
						10'd61	:	dt	<=	129	;
						10'd62	:	dt	<=	132	;
						10'd63	:	dt	<=	134	;
						10'd64	:	dt	<=	139	;
						10'd65	:	dt	<=	141	;
						10'd66	:	dt	<=	142	;
						10'd67	:	dt	<=	144	;
						10'd68	:	dt	<=	147	;
						10'd69	:	dt	<=	149	;
						10'd70	:	dt	<=	153	;
						10'd71	:	dt	<=	158	;
						10'd72	:	dt	<=	119	;
						10'd73	:	dt	<=	135	;
						10'd74	:	dt	<=	157	;
						10'd75	:	dt	<=	157	;
						10'd76	:	dt	<=	159	;
						10'd77	:	dt	<=	161	;
						10'd78	:	dt	<=	162	;
						10'd79	:	dt	<=	163	;
						10'd80	:	dt	<=	164	;
						10'd81	:	dt	<=	165	;
						10'd82	:	dt	<=	165	;
						10'd83	:	dt	<=	165	;
						10'd84	:	dt	<=	98	;
						10'd85	:	dt	<=	107	;
						10'd86	:	dt	<=	117	;
						10'd87	:	dt	<=	122	;
						10'd88	:	dt	<=	126	;
						10'd89	:	dt	<=	130	;
						10'd90	:	dt	<=	133	;
						10'd91	:	dt	<=	136	;
						10'd92	:	dt	<=	139	;
						10'd93	:	dt	<=	141	;
						10'd94	:	dt	<=	143	;
						10'd95	:	dt	<=	145	;
						10'd96	:	dt	<=	148	;
						10'd97	:	dt	<=	150	;
						10'd98	:	dt	<=	158	;
						10'd99	:	dt	<=	164	;
						10'd100	:	dt	<=	122	;
						10'd101	:	dt	<=	120	;
						10'd102	:	dt	<=	157	;
						10'd103	:	dt	<=	158	;
						10'd104	:	dt	<=	161	;
						10'd105	:	dt	<=	162	;
						10'd106	:	dt	<=	163	;
						10'd107	:	dt	<=	164	;
						10'd108	:	dt	<=	165	;
						10'd109	:	dt	<=	166	;
						10'd110	:	dt	<=	167	;
						10'd111	:	dt	<=	167	;
						10'd112	:	dt	<=	99	;
						10'd113	:	dt	<=	107	;
						10'd114	:	dt	<=	117	;
						10'd115	:	dt	<=	123	;
						10'd116	:	dt	<=	127	;
						10'd117	:	dt	<=	130	;
						10'd118	:	dt	<=	134	;
						10'd119	:	dt	<=	138	;
						10'd120	:	dt	<=	140	;
						10'd121	:	dt	<=	143	;
						10'd122	:	dt	<=	144	;
						10'd123	:	dt	<=	147	;
						10'd124	:	dt	<=	149	;
						10'd125	:	dt	<=	151	;
						10'd126	:	dt	<=	158	;
						10'd127	:	dt	<=	165	;
						10'd128	:	dt	<=	130	;
						10'd129	:	dt	<=	112	;
						10'd130	:	dt	<=	156	;
						10'd131	:	dt	<=	159	;
						10'd132	:	dt	<=	162	;
						10'd133	:	dt	<=	164	;
						10'd134	:	dt	<=	164	;
						10'd135	:	dt	<=	165	;
						10'd136	:	dt	<=	167	;
						10'd137	:	dt	<=	168	;
						10'd138	:	dt	<=	168	;
						10'd139	:	dt	<=	169	;
						10'd140	:	dt	<=	99	;
						10'd141	:	dt	<=	109	;
						10'd142	:	dt	<=	119	;
						10'd143	:	dt	<=	124	;
						10'd144	:	dt	<=	127	;
						10'd145	:	dt	<=	132	;
						10'd146	:	dt	<=	136	;
						10'd147	:	dt	<=	138	;
						10'd148	:	dt	<=	140	;
						10'd149	:	dt	<=	143	;
						10'd150	:	dt	<=	145	;
						10'd151	:	dt	<=	147	;
						10'd152	:	dt	<=	149	;
						10'd153	:	dt	<=	152	;
						10'd154	:	dt	<=	155	;
						10'd155	:	dt	<=	167	;
						10'd156	:	dt	<=	140	;
						10'd157	:	dt	<=	111	;
						10'd158	:	dt	<=	153	;
						10'd159	:	dt	<=	161	;
						10'd160	:	dt	<=	163	;
						10'd161	:	dt	<=	165	;
						10'd162	:	dt	<=	166	;
						10'd163	:	dt	<=	166	;
						10'd164	:	dt	<=	168	;
						10'd165	:	dt	<=	169	;
						10'd166	:	dt	<=	169	;
						10'd167	:	dt	<=	170	;
						10'd168	:	dt	<=	100	;
						10'd169	:	dt	<=	110	;
						10'd170	:	dt	<=	120	;
						10'd171	:	dt	<=	124	;
						10'd172	:	dt	<=	128	;
						10'd173	:	dt	<=	134	;
						10'd174	:	dt	<=	137	;
						10'd175	:	dt	<=	138	;
						10'd176	:	dt	<=	141	;
						10'd177	:	dt	<=	144	;
						10'd178	:	dt	<=	145	;
						10'd179	:	dt	<=	153	;
						10'd180	:	dt	<=	137	;
						10'd181	:	dt	<=	137	;
						10'd182	:	dt	<=	156	;
						10'd183	:	dt	<=	173	;
						10'd184	:	dt	<=	152	;
						10'd185	:	dt	<=	113	;
						10'd186	:	dt	<=	144	;
						10'd187	:	dt	<=	163	;
						10'd188	:	dt	<=	163	;
						10'd189	:	dt	<=	165	;
						10'd190	:	dt	<=	165	;
						10'd191	:	dt	<=	166	;
						10'd192	:	dt	<=	169	;
						10'd193	:	dt	<=	169	;
						10'd194	:	dt	<=	170	;
						10'd195	:	dt	<=	171	;
						10'd196	:	dt	<=	102	;
						10'd197	:	dt	<=	112	;
						10'd198	:	dt	<=	120	;
						10'd199	:	dt	<=	125	;
						10'd200	:	dt	<=	130	;
						10'd201	:	dt	<=	135	;
						10'd202	:	dt	<=	138	;
						10'd203	:	dt	<=	140	;
						10'd204	:	dt	<=	143	;
						10'd205	:	dt	<=	144	;
						10'd206	:	dt	<=	148	;
						10'd207	:	dt	<=	158	;
						10'd208	:	dt	<=	132	;
						10'd209	:	dt	<=	102	;
						10'd210	:	dt	<=	150	;
						10'd211	:	dt	<=	171	;
						10'd212	:	dt	<=	156	;
						10'd213	:	dt	<=	117	;
						10'd214	:	dt	<=	130	;
						10'd215	:	dt	<=	165	;
						10'd216	:	dt	<=	164	;
						10'd217	:	dt	<=	165	;
						10'd218	:	dt	<=	166	;
						10'd219	:	dt	<=	168	;
						10'd220	:	dt	<=	170	;
						10'd221	:	dt	<=	170	;
						10'd222	:	dt	<=	171	;
						10'd223	:	dt	<=	172	;
						10'd224	:	dt	<=	104	;
						10'd225	:	dt	<=	114	;
						10'd226	:	dt	<=	121	;
						10'd227	:	dt	<=	125	;
						10'd228	:	dt	<=	130	;
						10'd229	:	dt	<=	135	;
						10'd230	:	dt	<=	138	;
						10'd231	:	dt	<=	141	;
						10'd232	:	dt	<=	145	;
						10'd233	:	dt	<=	146	;
						10'd234	:	dt	<=	153	;
						10'd235	:	dt	<=	152	;
						10'd236	:	dt	<=	128	;
						10'd237	:	dt	<=	87	;
						10'd238	:	dt	<=	133	;
						10'd239	:	dt	<=	167	;
						10'd240	:	dt	<=	153	;
						10'd241	:	dt	<=	118	;
						10'd242	:	dt	<=	119	;
						10'd243	:	dt	<=	165	;
						10'd244	:	dt	<=	166	;
						10'd245	:	dt	<=	167	;
						10'd246	:	dt	<=	167	;
						10'd247	:	dt	<=	170	;
						10'd248	:	dt	<=	171	;
						10'd249	:	dt	<=	171	;
						10'd250	:	dt	<=	172	;
						10'd251	:	dt	<=	172	;
						10'd252	:	dt	<=	105	;
						10'd253	:	dt	<=	116	;
						10'd254	:	dt	<=	123	;
						10'd255	:	dt	<=	126	;
						10'd256	:	dt	<=	130	;
						10'd257	:	dt	<=	140	;
						10'd258	:	dt	<=	136	;
						10'd259	:	dt	<=	127	;
						10'd260	:	dt	<=	123	;
						10'd261	:	dt	<=	124	;
						10'd262	:	dt	<=	141	;
						10'd263	:	dt	<=	160	;
						10'd264	:	dt	<=	139	;
						10'd265	:	dt	<=	102	;
						10'd266	:	dt	<=	112	;
						10'd267	:	dt	<=	165	;
						10'd268	:	dt	<=	141	;
						10'd269	:	dt	<=	116	;
						10'd270	:	dt	<=	111	;
						10'd271	:	dt	<=	164	;
						10'd272	:	dt	<=	167	;
						10'd273	:	dt	<=	168	;
						10'd274	:	dt	<=	168	;
						10'd275	:	dt	<=	171	;
						10'd276	:	dt	<=	172	;
						10'd277	:	dt	<=	172	;
						10'd278	:	dt	<=	173	;
						10'd279	:	dt	<=	173	;
						10'd280	:	dt	<=	105	;
						10'd281	:	dt	<=	115	;
						10'd282	:	dt	<=	123	;
						10'd283	:	dt	<=	127	;
						10'd284	:	dt	<=	130	;
						10'd285	:	dt	<=	144	;
						10'd286	:	dt	<=	123	;
						10'd287	:	dt	<=	94	;
						10'd288	:	dt	<=	81	;
						10'd289	:	dt	<=	80	;
						10'd290	:	dt	<=	89	;
						10'd291	:	dt	<=	141	;
						10'd292	:	dt	<=	152	;
						10'd293	:	dt	<=	116	;
						10'd294	:	dt	<=	90	;
						10'd295	:	dt	<=	150	;
						10'd296	:	dt	<=	124	;
						10'd297	:	dt	<=	112	;
						10'd298	:	dt	<=	103	;
						10'd299	:	dt	<=	162	;
						10'd300	:	dt	<=	167	;
						10'd301	:	dt	<=	169	;
						10'd302	:	dt	<=	171	;
						10'd303	:	dt	<=	172	;
						10'd304	:	dt	<=	173	;
						10'd305	:	dt	<=	174	;
						10'd306	:	dt	<=	174	;
						10'd307	:	dt	<=	174	;
						10'd308	:	dt	<=	107	;
						10'd309	:	dt	<=	117	;
						10'd310	:	dt	<=	123	;
						10'd311	:	dt	<=	128	;
						10'd312	:	dt	<=	131	;
						10'd313	:	dt	<=	133	;
						10'd314	:	dt	<=	115	;
						10'd315	:	dt	<=	91	;
						10'd316	:	dt	<=	76	;
						10'd317	:	dt	<=	82	;
						10'd318	:	dt	<=	85	;
						10'd319	:	dt	<=	111	;
						10'd320	:	dt	<=	154	;
						10'd321	:	dt	<=	129	;
						10'd322	:	dt	<=	88	;
						10'd323	:	dt	<=	130	;
						10'd324	:	dt	<=	105	;
						10'd325	:	dt	<=	106	;
						10'd326	:	dt	<=	98	;
						10'd327	:	dt	<=	157	;
						10'd328	:	dt	<=	169	;
						10'd329	:	dt	<=	171	;
						10'd330	:	dt	<=	172	;
						10'd331	:	dt	<=	173	;
						10'd332	:	dt	<=	174	;
						10'd333	:	dt	<=	175	;
						10'd334	:	dt	<=	175	;
						10'd335	:	dt	<=	175	;
						10'd336	:	dt	<=	108	;
						10'd337	:	dt	<=	117	;
						10'd338	:	dt	<=	123	;
						10'd339	:	dt	<=	127	;
						10'd340	:	dt	<=	132	;
						10'd341	:	dt	<=	136	;
						10'd342	:	dt	<=	135	;
						10'd343	:	dt	<=	129	;
						10'd344	:	dt	<=	120	;
						10'd345	:	dt	<=	98	;
						10'd346	:	dt	<=	83	;
						10'd347	:	dt	<=	97	;
						10'd348	:	dt	<=	154	;
						10'd349	:	dt	<=	140	;
						10'd350	:	dt	<=	95	;
						10'd351	:	dt	<=	103	;
						10'd352	:	dt	<=	88	;
						10'd353	:	dt	<=	99	;
						10'd354	:	dt	<=	92	;
						10'd355	:	dt	<=	150	;
						10'd356	:	dt	<=	171	;
						10'd357	:	dt	<=	171	;
						10'd358	:	dt	<=	172	;
						10'd359	:	dt	<=	173	;
						10'd360	:	dt	<=	175	;
						10'd361	:	dt	<=	176	;
						10'd362	:	dt	<=	176	;
						10'd363	:	dt	<=	176	;
						10'd364	:	dt	<=	108	;
						10'd365	:	dt	<=	118	;
						10'd366	:	dt	<=	123	;
						10'd367	:	dt	<=	129	;
						10'd368	:	dt	<=	133	;
						10'd369	:	dt	<=	138	;
						10'd370	:	dt	<=	140	;
						10'd371	:	dt	<=	160	;
						10'd372	:	dt	<=	164	;
						10'd373	:	dt	<=	115	;
						10'd374	:	dt	<=	71	;
						10'd375	:	dt	<=	109	;
						10'd376	:	dt	<=	164	;
						10'd377	:	dt	<=	147	;
						10'd378	:	dt	<=	102	;
						10'd379	:	dt	<=	77	;
						10'd380	:	dt	<=	81	;
						10'd381	:	dt	<=	96	;
						10'd382	:	dt	<=	94	;
						10'd383	:	dt	<=	139	;
						10'd384	:	dt	<=	172	;
						10'd385	:	dt	<=	173	;
						10'd386	:	dt	<=	174	;
						10'd387	:	dt	<=	173	;
						10'd388	:	dt	<=	174	;
						10'd389	:	dt	<=	175	;
						10'd390	:	dt	<=	176	;
						10'd391	:	dt	<=	176	;
						10'd392	:	dt	<=	110	;
						10'd393	:	dt	<=	119	;
						10'd394	:	dt	<=	124	;
						10'd395	:	dt	<=	129	;
						10'd396	:	dt	<=	135	;
						10'd397	:	dt	<=	138	;
						10'd398	:	dt	<=	141	;
						10'd399	:	dt	<=	164	;
						10'd400	:	dt	<=	166	;
						10'd401	:	dt	<=	119	;
						10'd402	:	dt	<=	66	;
						10'd403	:	dt	<=	105	;
						10'd404	:	dt	<=	176	;
						10'd405	:	dt	<=	149	;
						10'd406	:	dt	<=	111	;
						10'd407	:	dt	<=	74	;
						10'd408	:	dt	<=	79	;
						10'd409	:	dt	<=	94	;
						10'd410	:	dt	<=	93	;
						10'd411	:	dt	<=	124	;
						10'd412	:	dt	<=	173	;
						10'd413	:	dt	<=	173	;
						10'd414	:	dt	<=	174	;
						10'd415	:	dt	<=	174	;
						10'd416	:	dt	<=	175	;
						10'd417	:	dt	<=	176	;
						10'd418	:	dt	<=	176	;
						10'd419	:	dt	<=	176	;
						10'd420	:	dt	<=	111	;
						10'd421	:	dt	<=	120	;
						10'd422	:	dt	<=	124	;
						10'd423	:	dt	<=	130	;
						10'd424	:	dt	<=	134	;
						10'd425	:	dt	<=	148	;
						10'd426	:	dt	<=	160	;
						10'd427	:	dt	<=	163	;
						10'd428	:	dt	<=	170	;
						10'd429	:	dt	<=	125	;
						10'd430	:	dt	<=	61	;
						10'd431	:	dt	<=	114	;
						10'd432	:	dt	<=	184	;
						10'd433	:	dt	<=	150	;
						10'd434	:	dt	<=	116	;
						10'd435	:	dt	<=	79	;
						10'd436	:	dt	<=	78	;
						10'd437	:	dt	<=	91	;
						10'd438	:	dt	<=	90	;
						10'd439	:	dt	<=	109	;
						10'd440	:	dt	<=	173	;
						10'd441	:	dt	<=	175	;
						10'd442	:	dt	<=	175	;
						10'd443	:	dt	<=	175	;
						10'd444	:	dt	<=	177	;
						10'd445	:	dt	<=	178	;
						10'd446	:	dt	<=	178	;
						10'd447	:	dt	<=	178	;
						10'd448	:	dt	<=	113	;
						10'd449	:	dt	<=	121	;
						10'd450	:	dt	<=	125	;
						10'd451	:	dt	<=	130	;
						10'd452	:	dt	<=	132	;
						10'd453	:	dt	<=	156	;
						10'd454	:	dt	<=	174	;
						10'd455	:	dt	<=	160	;
						10'd456	:	dt	<=	165	;
						10'd457	:	dt	<=	125	;
						10'd458	:	dt	<=	70	;
						10'd459	:	dt	<=	146	;
						10'd460	:	dt	<=	176	;
						10'd461	:	dt	<=	148	;
						10'd462	:	dt	<=	112	;
						10'd463	:	dt	<=	79	;
						10'd464	:	dt	<=	71	;
						10'd465	:	dt	<=	85	;
						10'd466	:	dt	<=	85	;
						10'd467	:	dt	<=	99	;
						10'd468	:	dt	<=	172	;
						10'd469	:	dt	<=	175	;
						10'd470	:	dt	<=	175	;
						10'd471	:	dt	<=	176	;
						10'd472	:	dt	<=	177	;
						10'd473	:	dt	<=	178	;
						10'd474	:	dt	<=	179	;
						10'd475	:	dt	<=	179	;
						10'd476	:	dt	<=	113	;
						10'd477	:	dt	<=	121	;
						10'd478	:	dt	<=	126	;
						10'd479	:	dt	<=	131	;
						10'd480	:	dt	<=	133	;
						10'd481	:	dt	<=	147	;
						10'd482	:	dt	<=	171	;
						10'd483	:	dt	<=	153	;
						10'd484	:	dt	<=	155	;
						10'd485	:	dt	<=	130	;
						10'd486	:	dt	<=	126	;
						10'd487	:	dt	<=	181	;
						10'd488	:	dt	<=	164	;
						10'd489	:	dt	<=	147	;
						10'd490	:	dt	<=	112	;
						10'd491	:	dt	<=	81	;
						10'd492	:	dt	<=	72	;
						10'd493	:	dt	<=	81	;
						10'd494	:	dt	<=	78	;
						10'd495	:	dt	<=	111	;
						10'd496	:	dt	<=	174	;
						10'd497	:	dt	<=	174	;
						10'd498	:	dt	<=	175	;
						10'd499	:	dt	<=	176	;
						10'd500	:	dt	<=	178	;
						10'd501	:	dt	<=	178	;
						10'd502	:	dt	<=	178	;
						10'd503	:	dt	<=	179	;
						10'd504	:	dt	<=	113	;
						10'd505	:	dt	<=	121	;
						10'd506	:	dt	<=	126	;
						10'd507	:	dt	<=	130	;
						10'd508	:	dt	<=	134	;
						10'd509	:	dt	<=	139	;
						10'd510	:	dt	<=	151	;
						10'd511	:	dt	<=	136	;
						10'd512	:	dt	<=	143	;
						10'd513	:	dt	<=	149	;
						10'd514	:	dt	<=	177	;
						10'd515	:	dt	<=	185	;
						10'd516	:	dt	<=	160	;
						10'd517	:	dt	<=	143	;
						10'd518	:	dt	<=	116	;
						10'd519	:	dt	<=	85	;
						10'd520	:	dt	<=	75	;
						10'd521	:	dt	<=	78	;
						10'd522	:	dt	<=	76	;
						10'd523	:	dt	<=	141	;
						10'd524	:	dt	<=	175	;
						10'd525	:	dt	<=	175	;
						10'd526	:	dt	<=	176	;
						10'd527	:	dt	<=	177	;
						10'd528	:	dt	<=	178	;
						10'd529	:	dt	<=	178	;
						10'd530	:	dt	<=	179	;
						10'd531	:	dt	<=	179	;
						10'd532	:	dt	<=	114	;
						10'd533	:	dt	<=	121	;
						10'd534	:	dt	<=	125	;
						10'd535	:	dt	<=	130	;
						10'd536	:	dt	<=	135	;
						10'd537	:	dt	<=	138	;
						10'd538	:	dt	<=	149	;
						10'd539	:	dt	<=	135	;
						10'd540	:	dt	<=	146	;
						10'd541	:	dt	<=	176	;
						10'd542	:	dt	<=	194	;
						10'd543	:	dt	<=	182	;
						10'd544	:	dt	<=	159	;
						10'd545	:	dt	<=	136	;
						10'd546	:	dt	<=	114	;
						10'd547	:	dt	<=	89	;
						10'd548	:	dt	<=	76	;
						10'd549	:	dt	<=	73	;
						10'd550	:	dt	<=	86	;
						10'd551	:	dt	<=	164	;
						10'd552	:	dt	<=	174	;
						10'd553	:	dt	<=	175	;
						10'd554	:	dt	<=	177	;
						10'd555	:	dt	<=	178	;
						10'd556	:	dt	<=	179	;
						10'd557	:	dt	<=	179	;
						10'd558	:	dt	<=	180	;
						10'd559	:	dt	<=	180	;
						10'd560	:	dt	<=	116	;
						10'd561	:	dt	<=	122	;
						10'd562	:	dt	<=	125	;
						10'd563	:	dt	<=	129	;
						10'd564	:	dt	<=	135	;
						10'd565	:	dt	<=	139	;
						10'd566	:	dt	<=	160	;
						10'd567	:	dt	<=	161	;
						10'd568	:	dt	<=	145	;
						10'd569	:	dt	<=	171	;
						10'd570	:	dt	<=	193	;
						10'd571	:	dt	<=	176	;
						10'd572	:	dt	<=	155	;
						10'd573	:	dt	<=	133	;
						10'd574	:	dt	<=	113	;
						10'd575	:	dt	<=	90	;
						10'd576	:	dt	<=	75	;
						10'd577	:	dt	<=	68	;
						10'd578	:	dt	<=	110	;
						10'd579	:	dt	<=	174	;
						10'd580	:	dt	<=	174	;
						10'd581	:	dt	<=	175	;
						10'd582	:	dt	<=	177	;
						10'd583	:	dt	<=	178	;
						10'd584	:	dt	<=	179	;
						10'd585	:	dt	<=	179	;
						10'd586	:	dt	<=	180	;
						10'd587	:	dt	<=	180	;
						10'd588	:	dt	<=	117	;
						10'd589	:	dt	<=	122	;
						10'd590	:	dt	<=	126	;
						10'd591	:	dt	<=	130	;
						10'd592	:	dt	<=	136	;
						10'd593	:	dt	<=	138	;
						10'd594	:	dt	<=	170	;
						10'd595	:	dt	<=	175	;
						10'd596	:	dt	<=	147	;
						10'd597	:	dt	<=	156	;
						10'd598	:	dt	<=	190	;
						10'd599	:	dt	<=	175	;
						10'd600	:	dt	<=	155	;
						10'd601	:	dt	<=	131	;
						10'd602	:	dt	<=	113	;
						10'd603	:	dt	<=	92	;
						10'd604	:	dt	<=	75	;
						10'd605	:	dt	<=	69	;
						10'd606	:	dt	<=	137	;
						10'd607	:	dt	<=	175	;
						10'd608	:	dt	<=	174	;
						10'd609	:	dt	<=	175	;
						10'd610	:	dt	<=	177	;
						10'd611	:	dt	<=	179	;
						10'd612	:	dt	<=	179	;
						10'd613	:	dt	<=	179	;
						10'd614	:	dt	<=	180	;
						10'd615	:	dt	<=	180	;
						10'd616	:	dt	<=	117	;
						10'd617	:	dt	<=	122	;
						10'd618	:	dt	<=	127	;
						10'd619	:	dt	<=	132	;
						10'd620	:	dt	<=	137	;
						10'd621	:	dt	<=	139	;
						10'd622	:	dt	<=	176	;
						10'd623	:	dt	<=	182	;
						10'd624	:	dt	<=	161	;
						10'd625	:	dt	<=	171	;
						10'd626	:	dt	<=	186	;
						10'd627	:	dt	<=	173	;
						10'd628	:	dt	<=	156	;
						10'd629	:	dt	<=	131	;
						10'd630	:	dt	<=	114	;
						10'd631	:	dt	<=	94	;
						10'd632	:	dt	<=	75	;
						10'd633	:	dt	<=	82	;
						10'd634	:	dt	<=	161	;
						10'd635	:	dt	<=	173	;
						10'd636	:	dt	<=	174	;
						10'd637	:	dt	<=	176	;
						10'd638	:	dt	<=	178	;
						10'd639	:	dt	<=	179	;
						10'd640	:	dt	<=	179	;
						10'd641	:	dt	<=	180	;
						10'd642	:	dt	<=	180	;
						10'd643	:	dt	<=	181	;
						10'd644	:	dt	<=	116	;
						10'd645	:	dt	<=	121	;
						10'd646	:	dt	<=	126	;
						10'd647	:	dt	<=	132	;
						10'd648	:	dt	<=	136	;
						10'd649	:	dt	<=	141	;
						10'd650	:	dt	<=	183	;
						10'd651	:	dt	<=	190	;
						10'd652	:	dt	<=	169	;
						10'd653	:	dt	<=	176	;
						10'd654	:	dt	<=	184	;
						10'd655	:	dt	<=	173	;
						10'd656	:	dt	<=	157	;
						10'd657	:	dt	<=	133	;
						10'd658	:	dt	<=	115	;
						10'd659	:	dt	<=	95	;
						10'd660	:	dt	<=	72	;
						10'd661	:	dt	<=	109	;
						10'd662	:	dt	<=	173	;
						10'd663	:	dt	<=	174	;
						10'd664	:	dt	<=	175	;
						10'd665	:	dt	<=	177	;
						10'd666	:	dt	<=	179	;
						10'd667	:	dt	<=	180	;
						10'd668	:	dt	<=	180	;
						10'd669	:	dt	<=	180	;
						10'd670	:	dt	<=	180	;
						10'd671	:	dt	<=	181	;
						10'd672	:	dt	<=	117	;
						10'd673	:	dt	<=	121	;
						10'd674	:	dt	<=	126	;
						10'd675	:	dt	<=	132	;
						10'd676	:	dt	<=	137	;
						10'd677	:	dt	<=	140	;
						10'd678	:	dt	<=	181	;
						10'd679	:	dt	<=	188	;
						10'd680	:	dt	<=	174	;
						10'd681	:	dt	<=	176	;
						10'd682	:	dt	<=	179	;
						10'd683	:	dt	<=	177	;
						10'd684	:	dt	<=	165	;
						10'd685	:	dt	<=	137	;
						10'd686	:	dt	<=	115	;
						10'd687	:	dt	<=	94	;
						10'd688	:	dt	<=	73	;
						10'd689	:	dt	<=	138	;
						10'd690	:	dt	<=	174	;
						10'd691	:	dt	<=	174	;
						10'd692	:	dt	<=	175	;
						10'd693	:	dt	<=	176	;
						10'd694	:	dt	<=	178	;
						10'd695	:	dt	<=	179	;
						10'd696	:	dt	<=	180	;
						10'd697	:	dt	<=	181	;
						10'd698	:	dt	<=	181	;
						10'd699	:	dt	<=	182	;
						10'd700	:	dt	<=	117	;
						10'd701	:	dt	<=	121	;
						10'd702	:	dt	<=	126	;
						10'd703	:	dt	<=	132	;
						10'd704	:	dt	<=	136	;
						10'd705	:	dt	<=	140	;
						10'd706	:	dt	<=	175	;
						10'd707	:	dt	<=	180	;
						10'd708	:	dt	<=	169	;
						10'd709	:	dt	<=	176	;
						10'd710	:	dt	<=	176	;
						10'd711	:	dt	<=	178	;
						10'd712	:	dt	<=	170	;
						10'd713	:	dt	<=	140	;
						10'd714	:	dt	<=	113	;
						10'd715	:	dt	<=	90	;
						10'd716	:	dt	<=	84	;
						10'd717	:	dt	<=	160	;
						10'd718	:	dt	<=	173	;
						10'd719	:	dt	<=	174	;
						10'd720	:	dt	<=	176	;
						10'd721	:	dt	<=	177	;
						10'd722	:	dt	<=	178	;
						10'd723	:	dt	<=	179	;
						10'd724	:	dt	<=	180	;
						10'd725	:	dt	<=	181	;
						10'd726	:	dt	<=	182	;
						10'd727	:	dt	<=	182	;
						10'd728	:	dt	<=	117	;
						10'd729	:	dt	<=	121	;
						10'd730	:	dt	<=	127	;
						10'd731	:	dt	<=	133	;
						10'd732	:	dt	<=	137	;
						10'd733	:	dt	<=	141	;
						10'd734	:	dt	<=	166	;
						10'd735	:	dt	<=	170	;
						10'd736	:	dt	<=	169	;
						10'd737	:	dt	<=	176	;
						10'd738	:	dt	<=	176	;
						10'd739	:	dt	<=	178	;
						10'd740	:	dt	<=	169	;
						10'd741	:	dt	<=	138	;
						10'd742	:	dt	<=	110	;
						10'd743	:	dt	<=	84	;
						10'd744	:	dt	<=	109	;
						10'd745	:	dt	<=	172	;
						10'd746	:	dt	<=	174	;
						10'd747	:	dt	<=	175	;
						10'd748	:	dt	<=	176	;
						10'd749	:	dt	<=	178	;
						10'd750	:	dt	<=	180	;
						10'd751	:	dt	<=	180	;
						10'd752	:	dt	<=	181	;
						10'd753	:	dt	<=	181	;
						10'd754	:	dt	<=	181	;
						10'd755	:	dt	<=	182	;
						10'd756	:	dt	<=	118	;
						10'd757	:	dt	<=	122	;
						10'd758	:	dt	<=	128	;
						10'd759	:	dt	<=	133	;
						10'd760	:	dt	<=	137	;
						10'd761	:	dt	<=	141	;
						10'd762	:	dt	<=	157	;
						10'd763	:	dt	<=	168	;
						10'd764	:	dt	<=	176	;
						10'd765	:	dt	<=	182	;
						10'd766	:	dt	<=	175	;
						10'd767	:	dt	<=	174	;
						10'd768	:	dt	<=	165	;
						10'd769	:	dt	<=	135	;
						10'd770	:	dt	<=	107	;
						10'd771	:	dt	<=	82	;
						10'd772	:	dt	<=	137	;
						10'd773	:	dt	<=	174	;
						10'd774	:	dt	<=	173	;
						10'd775	:	dt	<=	175	;
						10'd776	:	dt	<=	177	;
						10'd777	:	dt	<=	178	;
						10'd778	:	dt	<=	180	;
						10'd779	:	dt	<=	180	;
						10'd780	:	dt	<=	181	;
						10'd781	:	dt	<=	181	;
						10'd782	:	dt	<=	181	;
						10'd783	:	dt	<=	183	;
					endcase
				end
				5'd11	:	begin
					case (cnt)
						10'd0	:	dt	<=	84	;
						10'd1	:	dt	<=	89	;
						10'd2	:	dt	<=	95	;
						10'd3	:	dt	<=	101	;
						10'd4	:	dt	<=	104	;
						10'd5	:	dt	<=	108	;
						10'd6	:	dt	<=	112	;
						10'd7	:	dt	<=	116	;
						10'd8	:	dt	<=	118	;
						10'd9	:	dt	<=	120	;
						10'd10	:	dt	<=	122	;
						10'd11	:	dt	<=	122	;
						10'd12	:	dt	<=	124	;
						10'd13	:	dt	<=	128	;
						10'd14	:	dt	<=	127	;
						10'd15	:	dt	<=	127	;
						10'd16	:	dt	<=	127	;
						10'd17	:	dt	<=	127	;
						10'd18	:	dt	<=	127	;
						10'd19	:	dt	<=	127	;
						10'd20	:	dt	<=	127	;
						10'd21	:	dt	<=	126	;
						10'd22	:	dt	<=	124	;
						10'd23	:	dt	<=	128	;
						10'd24	:	dt	<=	93	;
						10'd25	:	dt	<=	70	;
						10'd26	:	dt	<=	110	;
						10'd27	:	dt	<=	148	;
						10'd28	:	dt	<=	87	;
						10'd29	:	dt	<=	91	;
						10'd30	:	dt	<=	96	;
						10'd31	:	dt	<=	102	;
						10'd32	:	dt	<=	106	;
						10'd33	:	dt	<=	110	;
						10'd34	:	dt	<=	113	;
						10'd35	:	dt	<=	116	;
						10'd36	:	dt	<=	119	;
						10'd37	:	dt	<=	121	;
						10'd38	:	dt	<=	123	;
						10'd39	:	dt	<=	122	;
						10'd40	:	dt	<=	140	;
						10'd41	:	dt	<=	113	;
						10'd42	:	dt	<=	126	;
						10'd43	:	dt	<=	126	;
						10'd44	:	dt	<=	127	;
						10'd45	:	dt	<=	127	;
						10'd46	:	dt	<=	126	;
						10'd47	:	dt	<=	126	;
						10'd48	:	dt	<=	126	;
						10'd49	:	dt	<=	124	;
						10'd50	:	dt	<=	122	;
						10'd51	:	dt	<=	127	;
						10'd52	:	dt	<=	100	;
						10'd53	:	dt	<=	86	;
						10'd54	:	dt	<=	111	;
						10'd55	:	dt	<=	152	;
						10'd56	:	dt	<=	90	;
						10'd57	:	dt	<=	95	;
						10'd58	:	dt	<=	100	;
						10'd59	:	dt	<=	106	;
						10'd60	:	dt	<=	109	;
						10'd61	:	dt	<=	113	;
						10'd62	:	dt	<=	116	;
						10'd63	:	dt	<=	120	;
						10'd64	:	dt	<=	122	;
						10'd65	:	dt	<=	124	;
						10'd66	:	dt	<=	126	;
						10'd67	:	dt	<=	122	;
						10'd68	:	dt	<=	159	;
						10'd69	:	dt	<=	94	;
						10'd70	:	dt	<=	109	;
						10'd71	:	dt	<=	132	;
						10'd72	:	dt	<=	126	;
						10'd73	:	dt	<=	128	;
						10'd74	:	dt	<=	127	;
						10'd75	:	dt	<=	127	;
						10'd76	:	dt	<=	126	;
						10'd77	:	dt	<=	124	;
						10'd78	:	dt	<=	124	;
						10'd79	:	dt	<=	121	;
						10'd80	:	dt	<=	112	;
						10'd81	:	dt	<=	150	;
						10'd82	:	dt	<=	144	;
						10'd83	:	dt	<=	147	;
						10'd84	:	dt	<=	93	;
						10'd85	:	dt	<=	98	;
						10'd86	:	dt	<=	105	;
						10'd87	:	dt	<=	110	;
						10'd88	:	dt	<=	115	;
						10'd89	:	dt	<=	118	;
						10'd90	:	dt	<=	122	;
						10'd91	:	dt	<=	125	;
						10'd92	:	dt	<=	127	;
						10'd93	:	dt	<=	128	;
						10'd94	:	dt	<=	130	;
						10'd95	:	dt	<=	127	;
						10'd96	:	dt	<=	172	;
						10'd97	:	dt	<=	101	;
						10'd98	:	dt	<=	87	;
						10'd99	:	dt	<=	138	;
						10'd100	:	dt	<=	128	;
						10'd101	:	dt	<=	129	;
						10'd102	:	dt	<=	129	;
						10'd103	:	dt	<=	128	;
						10'd104	:	dt	<=	127	;
						10'd105	:	dt	<=	126	;
						10'd106	:	dt	<=	125	;
						10'd107	:	dt	<=	119	;
						10'd108	:	dt	<=	137	;
						10'd109	:	dt	<=	122	;
						10'd110	:	dt	<=	145	;
						10'd111	:	dt	<=	148	;
						10'd112	:	dt	<=	98	;
						10'd113	:	dt	<=	102	;
						10'd114	:	dt	<=	109	;
						10'd115	:	dt	<=	115	;
						10'd116	:	dt	<=	119	;
						10'd117	:	dt	<=	124	;
						10'd118	:	dt	<=	127	;
						10'd119	:	dt	<=	131	;
						10'd120	:	dt	<=	133	;
						10'd121	:	dt	<=	134	;
						10'd122	:	dt	<=	135	;
						10'd123	:	dt	<=	134	;
						10'd124	:	dt	<=	175	;
						10'd125	:	dt	<=	97	;
						10'd126	:	dt	<=	78	;
						10'd127	:	dt	<=	141	;
						10'd128	:	dt	<=	134	;
						10'd129	:	dt	<=	133	;
						10'd130	:	dt	<=	133	;
						10'd131	:	dt	<=	132	;
						10'd132	:	dt	<=	131	;
						10'd133	:	dt	<=	130	;
						10'd134	:	dt	<=	129	;
						10'd135	:	dt	<=	128	;
						10'd136	:	dt	<=	131	;
						10'd137	:	dt	<=	102	;
						10'd138	:	dt	<=	154	;
						10'd139	:	dt	<=	148	;
						10'd140	:	dt	<=	101	;
						10'd141	:	dt	<=	107	;
						10'd142	:	dt	<=	116	;
						10'd143	:	dt	<=	121	;
						10'd144	:	dt	<=	124	;
						10'd145	:	dt	<=	129	;
						10'd146	:	dt	<=	133	;
						10'd147	:	dt	<=	136	;
						10'd148	:	dt	<=	139	;
						10'd149	:	dt	<=	140	;
						10'd150	:	dt	<=	141	;
						10'd151	:	dt	<=	141	;
						10'd152	:	dt	<=	174	;
						10'd153	:	dt	<=	89	;
						10'd154	:	dt	<=	84	;
						10'd155	:	dt	<=	147	;
						10'd156	:	dt	<=	138	;
						10'd157	:	dt	<=	140	;
						10'd158	:	dt	<=	139	;
						10'd159	:	dt	<=	138	;
						10'd160	:	dt	<=	136	;
						10'd161	:	dt	<=	135	;
						10'd162	:	dt	<=	134	;
						10'd163	:	dt	<=	130	;
						10'd164	:	dt	<=	133	;
						10'd165	:	dt	<=	149	;
						10'd166	:	dt	<=	143	;
						10'd167	:	dt	<=	148	;
						10'd168	:	dt	<=	104	;
						10'd169	:	dt	<=	110	;
						10'd170	:	dt	<=	120	;
						10'd171	:	dt	<=	127	;
						10'd172	:	dt	<=	131	;
						10'd173	:	dt	<=	134	;
						10'd174	:	dt	<=	138	;
						10'd175	:	dt	<=	142	;
						10'd176	:	dt	<=	145	;
						10'd177	:	dt	<=	147	;
						10'd178	:	dt	<=	146	;
						10'd179	:	dt	<=	151	;
						10'd180	:	dt	<=	181	;
						10'd181	:	dt	<=	86	;
						10'd182	:	dt	<=	91	;
						10'd183	:	dt	<=	154	;
						10'd184	:	dt	<=	144	;
						10'd185	:	dt	<=	145	;
						10'd186	:	dt	<=	144	;
						10'd187	:	dt	<=	144	;
						10'd188	:	dt	<=	142	;
						10'd189	:	dt	<=	140	;
						10'd190	:	dt	<=	137	;
						10'd191	:	dt	<=	135	;
						10'd192	:	dt	<=	136	;
						10'd193	:	dt	<=	121	;
						10'd194	:	dt	<=	109	;
						10'd195	:	dt	<=	150	;
						10'd196	:	dt	<=	106	;
						10'd197	:	dt	<=	114	;
						10'd198	:	dt	<=	124	;
						10'd199	:	dt	<=	132	;
						10'd200	:	dt	<=	136	;
						10'd201	:	dt	<=	140	;
						10'd202	:	dt	<=	144	;
						10'd203	:	dt	<=	147	;
						10'd204	:	dt	<=	150	;
						10'd205	:	dt	<=	153	;
						10'd206	:	dt	<=	148	;
						10'd207	:	dt	<=	171	;
						10'd208	:	dt	<=	184	;
						10'd209	:	dt	<=	64	;
						10'd210	:	dt	<=	108	;
						10'd211	:	dt	<=	160	;
						10'd212	:	dt	<=	149	;
						10'd213	:	dt	<=	149	;
						10'd214	:	dt	<=	149	;
						10'd215	:	dt	<=	148	;
						10'd216	:	dt	<=	147	;
						10'd217	:	dt	<=	145	;
						10'd218	:	dt	<=	143	;
						10'd219	:	dt	<=	140	;
						10'd220	:	dt	<=	139	;
						10'd221	:	dt	<=	130	;
						10'd222	:	dt	<=	130	;
						10'd223	:	dt	<=	148	;
						10'd224	:	dt	<=	110	;
						10'd225	:	dt	<=	118	;
						10'd226	:	dt	<=	130	;
						10'd227	:	dt	<=	136	;
						10'd228	:	dt	<=	140	;
						10'd229	:	dt	<=	145	;
						10'd230	:	dt	<=	150	;
						10'd231	:	dt	<=	154	;
						10'd232	:	dt	<=	155	;
						10'd233	:	dt	<=	158	;
						10'd234	:	dt	<=	152	;
						10'd235	:	dt	<=	178	;
						10'd236	:	dt	<=	166	;
						10'd237	:	dt	<=	64	;
						10'd238	:	dt	<=	126	;
						10'd239	:	dt	<=	165	;
						10'd240	:	dt	<=	155	;
						10'd241	:	dt	<=	155	;
						10'd242	:	dt	<=	155	;
						10'd243	:	dt	<=	153	;
						10'd244	:	dt	<=	152	;
						10'd245	:	dt	<=	150	;
						10'd246	:	dt	<=	148	;
						10'd247	:	dt	<=	145	;
						10'd248	:	dt	<=	144	;
						10'd249	:	dt	<=	140	;
						10'd250	:	dt	<=	144	;
						10'd251	:	dt	<=	154	;
						10'd252	:	dt	<=	112	;
						10'd253	:	dt	<=	122	;
						10'd254	:	dt	<=	133	;
						10'd255	:	dt	<=	140	;
						10'd256	:	dt	<=	145	;
						10'd257	:	dt	<=	149	;
						10'd258	:	dt	<=	154	;
						10'd259	:	dt	<=	158	;
						10'd260	:	dt	<=	160	;
						10'd261	:	dt	<=	159	;
						10'd262	:	dt	<=	174	;
						10'd263	:	dt	<=	177	;
						10'd264	:	dt	<=	91	;
						10'd265	:	dt	<=	56	;
						10'd266	:	dt	<=	135	;
						10'd267	:	dt	<=	168	;
						10'd268	:	dt	<=	159	;
						10'd269	:	dt	<=	159	;
						10'd270	:	dt	<=	158	;
						10'd271	:	dt	<=	158	;
						10'd272	:	dt	<=	157	;
						10'd273	:	dt	<=	155	;
						10'd274	:	dt	<=	152	;
						10'd275	:	dt	<=	151	;
						10'd276	:	dt	<=	148	;
						10'd277	:	dt	<=	144	;
						10'd278	:	dt	<=	147	;
						10'd279	:	dt	<=	164	;
						10'd280	:	dt	<=	116	;
						10'd281	:	dt	<=	125	;
						10'd282	:	dt	<=	137	;
						10'd283	:	dt	<=	144	;
						10'd284	:	dt	<=	149	;
						10'd285	:	dt	<=	154	;
						10'd286	:	dt	<=	158	;
						10'd287	:	dt	<=	161	;
						10'd288	:	dt	<=	161	;
						10'd289	:	dt	<=	164	;
						10'd290	:	dt	<=	163	;
						10'd291	:	dt	<=	167	;
						10'd292	:	dt	<=	97	;
						10'd293	:	dt	<=	56	;
						10'd294	:	dt	<=	144	;
						10'd295	:	dt	<=	170	;
						10'd296	:	dt	<=	164	;
						10'd297	:	dt	<=	164	;
						10'd298	:	dt	<=	164	;
						10'd299	:	dt	<=	163	;
						10'd300	:	dt	<=	162	;
						10'd301	:	dt	<=	159	;
						10'd302	:	dt	<=	157	;
						10'd303	:	dt	<=	155	;
						10'd304	:	dt	<=	152	;
						10'd305	:	dt	<=	148	;
						10'd306	:	dt	<=	148	;
						10'd307	:	dt	<=	165	;
						10'd308	:	dt	<=	119	;
						10'd309	:	dt	<=	129	;
						10'd310	:	dt	<=	140	;
						10'd311	:	dt	<=	147	;
						10'd312	:	dt	<=	151	;
						10'd313	:	dt	<=	157	;
						10'd314	:	dt	<=	161	;
						10'd315	:	dt	<=	167	;
						10'd316	:	dt	<=	186	;
						10'd317	:	dt	<=	182	;
						10'd318	:	dt	<=	84	;
						10'd319	:	dt	<=	82	;
						10'd320	:	dt	<=	118	;
						10'd321	:	dt	<=	69	;
						10'd322	:	dt	<=	149	;
						10'd323	:	dt	<=	173	;
						10'd324	:	dt	<=	167	;
						10'd325	:	dt	<=	168	;
						10'd326	:	dt	<=	168	;
						10'd327	:	dt	<=	167	;
						10'd328	:	dt	<=	166	;
						10'd329	:	dt	<=	163	;
						10'd330	:	dt	<=	161	;
						10'd331	:	dt	<=	160	;
						10'd332	:	dt	<=	156	;
						10'd333	:	dt	<=	154	;
						10'd334	:	dt	<=	156	;
						10'd335	:	dt	<=	165	;
						10'd336	:	dt	<=	122	;
						10'd337	:	dt	<=	132	;
						10'd338	:	dt	<=	143	;
						10'd339	:	dt	<=	150	;
						10'd340	:	dt	<=	155	;
						10'd341	:	dt	<=	158	;
						10'd342	:	dt	<=	164	;
						10'd343	:	dt	<=	153	;
						10'd344	:	dt	<=	174	;
						10'd345	:	dt	<=	169	;
						10'd346	:	dt	<=	95	;
						10'd347	:	dt	<=	59	;
						10'd348	:	dt	<=	111	;
						10'd349	:	dt	<=	83	;
						10'd350	:	dt	<=	133	;
						10'd351	:	dt	<=	180	;
						10'd352	:	dt	<=	169	;
						10'd353	:	dt	<=	170	;
						10'd354	:	dt	<=	171	;
						10'd355	:	dt	<=	170	;
						10'd356	:	dt	<=	168	;
						10'd357	:	dt	<=	166	;
						10'd358	:	dt	<=	164	;
						10'd359	:	dt	<=	162	;
						10'd360	:	dt	<=	161	;
						10'd361	:	dt	<=	149	;
						10'd362	:	dt	<=	136	;
						10'd363	:	dt	<=	168	;
						10'd364	:	dt	<=	123	;
						10'd365	:	dt	<=	134	;
						10'd366	:	dt	<=	146	;
						10'd367	:	dt	<=	154	;
						10'd368	:	dt	<=	156	;
						10'd369	:	dt	<=	163	;
						10'd370	:	dt	<=	189	;
						10'd371	:	dt	<=	136	;
						10'd372	:	dt	<=	70	;
						10'd373	:	dt	<=	106	;
						10'd374	:	dt	<=	131	;
						10'd375	:	dt	<=	74	;
						10'd376	:	dt	<=	89	;
						10'd377	:	dt	<=	83	;
						10'd378	:	dt	<=	112	;
						10'd379	:	dt	<=	184	;
						10'd380	:	dt	<=	172	;
						10'd381	:	dt	<=	174	;
						10'd382	:	dt	<=	174	;
						10'd383	:	dt	<=	173	;
						10'd384	:	dt	<=	173	;
						10'd385	:	dt	<=	171	;
						10'd386	:	dt	<=	170	;
						10'd387	:	dt	<=	166	;
						10'd388	:	dt	<=	176	;
						10'd389	:	dt	<=	94	;
						10'd390	:	dt	<=	66	;
						10'd391	:	dt	<=	173	;
						10'd392	:	dt	<=	126	;
						10'd393	:	dt	<=	137	;
						10'd394	:	dt	<=	149	;
						10'd395	:	dt	<=	153	;
						10'd396	:	dt	<=	167	;
						10'd397	:	dt	<=	190	;
						10'd398	:	dt	<=	178	;
						10'd399	:	dt	<=	153	;
						10'd400	:	dt	<=	111	;
						10'd401	:	dt	<=	66	;
						10'd402	:	dt	<=	115	;
						10'd403	:	dt	<=	91	;
						10'd404	:	dt	<=	65	;
						10'd405	:	dt	<=	89	;
						10'd406	:	dt	<=	83	;
						10'd407	:	dt	<=	181	;
						10'd408	:	dt	<=	176	;
						10'd409	:	dt	<=	178	;
						10'd410	:	dt	<=	178	;
						10'd411	:	dt	<=	174	;
						10'd412	:	dt	<=	169	;
						10'd413	:	dt	<=	157	;
						10'd414	:	dt	<=	142	;
						10'd415	:	dt	<=	140	;
						10'd416	:	dt	<=	136	;
						10'd417	:	dt	<=	58	;
						10'd418	:	dt	<=	40	;
						10'd419	:	dt	<=	72	;
						10'd420	:	dt	<=	128	;
						10'd421	:	dt	<=	140	;
						10'd422	:	dt	<=	149	;
						10'd423	:	dt	<=	166	;
						10'd424	:	dt	<=	191	;
						10'd425	:	dt	<=	153	;
						10'd426	:	dt	<=	110	;
						10'd427	:	dt	<=	137	;
						10'd428	:	dt	<=	152	;
						10'd429	:	dt	<=	85	;
						10'd430	:	dt	<=	69	;
						10'd431	:	dt	<=	81	;
						10'd432	:	dt	<=	57	;
						10'd433	:	dt	<=	104	;
						10'd434	:	dt	<=	77	;
						10'd435	:	dt	<=	165	;
						10'd436	:	dt	<=	187	;
						10'd437	:	dt	<=	179	;
						10'd438	:	dt	<=	171	;
						10'd439	:	dt	<=	164	;
						10'd440	:	dt	<=	169	;
						10'd441	:	dt	<=	149	;
						10'd442	:	dt	<=	127	;
						10'd443	:	dt	<=	125	;
						10'd444	:	dt	<=	104	;
						10'd445	:	dt	<=	60	;
						10'd446	:	dt	<=	47	;
						10'd447	:	dt	<=	37	;
						10'd448	:	dt	<=	129	;
						10'd449	:	dt	<=	143	;
						10'd450	:	dt	<=	150	;
						10'd451	:	dt	<=	188	;
						10'd452	:	dt	<=	176	;
						10'd453	:	dt	<=	116	;
						10'd454	:	dt	<=	79	;
						10'd455	:	dt	<=	70	;
						10'd456	:	dt	<=	140	;
						10'd457	:	dt	<=	93	;
						10'd458	:	dt	<=	54	;
						10'd459	:	dt	<=	74	;
						10'd460	:	dt	<=	47	;
						10'd461	:	dt	<=	120	;
						10'd462	:	dt	<=	116	;
						10'd463	:	dt	<=	120	;
						10'd464	:	dt	<=	172	;
						10'd465	:	dt	<=	170	;
						10'd466	:	dt	<=	176	;
						10'd467	:	dt	<=	175	;
						10'd468	:	dt	<=	165	;
						10'd469	:	dt	<=	139	;
						10'd470	:	dt	<=	113	;
						10'd471	:	dt	<=	93	;
						10'd472	:	dt	<=	73	;
						10'd473	:	dt	<=	51	;
						10'd474	:	dt	<=	43	;
						10'd475	:	dt	<=	43	;
						10'd476	:	dt	<=	132	;
						10'd477	:	dt	<=	143	;
						10'd478	:	dt	<=	153	;
						10'd479	:	dt	<=	185	;
						10'd480	:	dt	<=	156	;
						10'd481	:	dt	<=	100	;
						10'd482	:	dt	<=	73	;
						10'd483	:	dt	<=	40	;
						10'd484	:	dt	<=	110	;
						10'd485	:	dt	<=	100	;
						10'd486	:	dt	<=	57	;
						10'd487	:	dt	<=	86	;
						10'd488	:	dt	<=	40	;
						10'd489	:	dt	<=	84	;
						10'd490	:	dt	<=	126	;
						10'd491	:	dt	<=	71	;
						10'd492	:	dt	<=	132	;
						10'd493	:	dt	<=	176	;
						10'd494	:	dt	<=	178	;
						10'd495	:	dt	<=	153	;
						10'd496	:	dt	<=	114	;
						10'd497	:	dt	<=	83	;
						10'd498	:	dt	<=	48	;
						10'd499	:	dt	<=	30	;
						10'd500	:	dt	<=	40	;
						10'd501	:	dt	<=	36	;
						10'd502	:	dt	<=	39	;
						10'd503	:	dt	<=	42	;
						10'd504	:	dt	<=	133	;
						10'd505	:	dt	<=	145	;
						10'd506	:	dt	<=	152	;
						10'd507	:	dt	<=	175	;
						10'd508	:	dt	<=	139	;
						10'd509	:	dt	<=	89	;
						10'd510	:	dt	<=	67	;
						10'd511	:	dt	<=	47	;
						10'd512	:	dt	<=	80	;
						10'd513	:	dt	<=	109	;
						10'd514	:	dt	<=	65	;
						10'd515	:	dt	<=	100	;
						10'd516	:	dt	<=	62	;
						10'd517	:	dt	<=	90	;
						10'd518	:	dt	<=	117	;
						10'd519	:	dt	<=	105	;
						10'd520	:	dt	<=	146	;
						10'd521	:	dt	<=	159	;
						10'd522	:	dt	<=	132	;
						10'd523	:	dt	<=	85	;
						10'd524	:	dt	<=	57	;
						10'd525	:	dt	<=	37	;
						10'd526	:	dt	<=	27	;
						10'd527	:	dt	<=	30	;
						10'd528	:	dt	<=	30	;
						10'd529	:	dt	<=	30	;
						10'd530	:	dt	<=	32	;
						10'd531	:	dt	<=	40	;
						10'd532	:	dt	<=	135	;
						10'd533	:	dt	<=	147	;
						10'd534	:	dt	<=	153	;
						10'd535	:	dt	<=	175	;
						10'd536	:	dt	<=	157	;
						10'd537	:	dt	<=	108	;
						10'd538	:	dt	<=	80	;
						10'd539	:	dt	<=	62	;
						10'd540	:	dt	<=	61	;
						10'd541	:	dt	<=	89	;
						10'd542	:	dt	<=	84	;
						10'd543	:	dt	<=	109	;
						10'd544	:	dt	<=	90	;
						10'd545	:	dt	<=	155	;
						10'd546	:	dt	<=	130	;
						10'd547	:	dt	<=	101	;
						10'd548	:	dt	<=	121	;
						10'd549	:	dt	<=	104	;
						10'd550	:	dt	<=	62	;
						10'd551	:	dt	<=	28	;
						10'd552	:	dt	<=	36	;
						10'd553	:	dt	<=	42	;
						10'd554	:	dt	<=	27	;
						10'd555	:	dt	<=	25	;
						10'd556	:	dt	<=	27	;
						10'd557	:	dt	<=	28	;
						10'd558	:	dt	<=	37	;
						10'd559	:	dt	<=	10	;
						10'd560	:	dt	<=	134	;
						10'd561	:	dt	<=	147	;
						10'd562	:	dt	<=	154	;
						10'd563	:	dt	<=	180	;
						10'd564	:	dt	<=	162	;
						10'd565	:	dt	<=	115	;
						10'd566	:	dt	<=	92	;
						10'd567	:	dt	<=	70	;
						10'd568	:	dt	<=	68	;
						10'd569	:	dt	<=	80	;
						10'd570	:	dt	<=	122	;
						10'd571	:	dt	<=	155	;
						10'd572	:	dt	<=	160	;
						10'd573	:	dt	<=	156	;
						10'd574	:	dt	<=	115	;
						10'd575	:	dt	<=	89	;
						10'd576	:	dt	<=	87	;
						10'd577	:	dt	<=	32	;
						10'd578	:	dt	<=	26	;
						10'd579	:	dt	<=	30	;
						10'd580	:	dt	<=	22	;
						10'd581	:	dt	<=	38	;
						10'd582	:	dt	<=	38	;
						10'd583	:	dt	<=	20	;
						10'd584	:	dt	<=	19	;
						10'd585	:	dt	<=	26	;
						10'd586	:	dt	<=	26	;
						10'd587	:	dt	<=	5	;
						10'd588	:	dt	<=	134	;
						10'd589	:	dt	<=	147	;
						10'd590	:	dt	<=	154	;
						10'd591	:	dt	<=	181	;
						10'd592	:	dt	<=	167	;
						10'd593	:	dt	<=	132	;
						10'd594	:	dt	<=	104	;
						10'd595	:	dt	<=	75	;
						10'd596	:	dt	<=	82	;
						10'd597	:	dt	<=	91	;
						10'd598	:	dt	<=	160	;
						10'd599	:	dt	<=	188	;
						10'd600	:	dt	<=	175	;
						10'd601	:	dt	<=	136	;
						10'd602	:	dt	<=	97	;
						10'd603	:	dt	<=	77	;
						10'd604	:	dt	<=	41	;
						10'd605	:	dt	<=	26	;
						10'd606	:	dt	<=	14	;
						10'd607	:	dt	<=	36	;
						10'd608	:	dt	<=	23	;
						10'd609	:	dt	<=	21	;
						10'd610	:	dt	<=	38	;
						10'd611	:	dt	<=	32	;
						10'd612	:	dt	<=	16	;
						10'd613	:	dt	<=	16	;
						10'd614	:	dt	<=	16	;
						10'd615	:	dt	<=	18	;
						10'd616	:	dt	<=	134	;
						10'd617	:	dt	<=	147	;
						10'd618	:	dt	<=	154	;
						10'd619	:	dt	<=	177	;
						10'd620	:	dt	<=	167	;
						10'd621	:	dt	<=	141	;
						10'd622	:	dt	<=	107	;
						10'd623	:	dt	<=	84	;
						10'd624	:	dt	<=	92	;
						10'd625	:	dt	<=	99	;
						10'd626	:	dt	<=	166	;
						10'd627	:	dt	<=	174	;
						10'd628	:	dt	<=	146	;
						10'd629	:	dt	<=	114	;
						10'd630	:	dt	<=	88	;
						10'd631	:	dt	<=	46	;
						10'd632	:	dt	<=	3	;
						10'd633	:	dt	<=	35	;
						10'd634	:	dt	<=	21	;
						10'd635	:	dt	<=	17	;
						10'd636	:	dt	<=	33	;
						10'd637	:	dt	<=	22	;
						10'd638	:	dt	<=	24	;
						10'd639	:	dt	<=	33	;
						10'd640	:	dt	<=	25	;
						10'd641	:	dt	<=	14	;
						10'd642	:	dt	<=	16	;
						10'd643	:	dt	<=	16	;
						10'd644	:	dt	<=	138	;
						10'd645	:	dt	<=	151	;
						10'd646	:	dt	<=	162	;
						10'd647	:	dt	<=	171	;
						10'd648	:	dt	<=	162	;
						10'd649	:	dt	<=	149	;
						10'd650	:	dt	<=	114	;
						10'd651	:	dt	<=	99	;
						10'd652	:	dt	<=	98	;
						10'd653	:	dt	<=	102	;
						10'd654	:	dt	<=	150	;
						10'd655	:	dt	<=	164	;
						10'd656	:	dt	<=	130	;
						10'd657	:	dt	<=	96	;
						10'd658	:	dt	<=	77	;
						10'd659	:	dt	<=	43	;
						10'd660	:	dt	<=	0	;
						10'd661	:	dt	<=	16	;
						10'd662	:	dt	<=	36	;
						10'd663	:	dt	<=	15	;
						10'd664	:	dt	<=	24	;
						10'd665	:	dt	<=	31	;
						10'd666	:	dt	<=	19	;
						10'd667	:	dt	<=	20	;
						10'd668	:	dt	<=	29	;
						10'd669	:	dt	<=	16	;
						10'd670	:	dt	<=	14	;
						10'd671	:	dt	<=	15	;
						10'd672	:	dt	<=	108	;
						10'd673	:	dt	<=	116	;
						10'd674	:	dt	<=	121	;
						10'd675	:	dt	<=	134	;
						10'd676	:	dt	<=	163	;
						10'd677	:	dt	<=	152	;
						10'd678	:	dt	<=	120	;
						10'd679	:	dt	<=	113	;
						10'd680	:	dt	<=	99	;
						10'd681	:	dt	<=	101	;
						10'd682	:	dt	<=	134	;
						10'd683	:	dt	<=	151	;
						10'd684	:	dt	<=	123	;
						10'd685	:	dt	<=	91	;
						10'd686	:	dt	<=	54	;
						10'd687	:	dt	<=	34	;
						10'd688	:	dt	<=	14	;
						10'd689	:	dt	<=	1	;
						10'd690	:	dt	<=	33	;
						10'd691	:	dt	<=	29	;
						10'd692	:	dt	<=	15	;
						10'd693	:	dt	<=	25	;
						10'd694	:	dt	<=	27	;
						10'd695	:	dt	<=	15	;
						10'd696	:	dt	<=	20	;
						10'd697	:	dt	<=	23	;
						10'd698	:	dt	<=	8	;
						10'd699	:	dt	<=	15	;
						10'd700	:	dt	<=	84	;
						10'd701	:	dt	<=	84	;
						10'd702	:	dt	<=	79	;
						10'd703	:	dt	<=	96	;
						10'd704	:	dt	<=	162	;
						10'd705	:	dt	<=	148	;
						10'd706	:	dt	<=	127	;
						10'd707	:	dt	<=	119	;
						10'd708	:	dt	<=	99	;
						10'd709	:	dt	<=	90	;
						10'd710	:	dt	<=	123	;
						10'd711	:	dt	<=	125	;
						10'd712	:	dt	<=	101	;
						10'd713	:	dt	<=	67	;
						10'd714	:	dt	<=	14	;
						10'd715	:	dt	<=	24	;
						10'd716	:	dt	<=	28	;
						10'd717	:	dt	<=	0	;
						10'd718	:	dt	<=	19	;
						10'd719	:	dt	<=	33	;
						10'd720	:	dt	<=	23	;
						10'd721	:	dt	<=	20	;
						10'd722	:	dt	<=	23	;
						10'd723	:	dt	<=	18	;
						10'd724	:	dt	<=	12	;
						10'd725	:	dt	<=	22	;
						10'd726	:	dt	<=	12	;
						10'd727	:	dt	<=	5	;
						10'd728	:	dt	<=	90	;
						10'd729	:	dt	<=	90	;
						10'd730	:	dt	<=	87	;
						10'd731	:	dt	<=	102	;
						10'd732	:	dt	<=	167	;
						10'd733	:	dt	<=	152	;
						10'd734	:	dt	<=	132	;
						10'd735	:	dt	<=	118	;
						10'd736	:	dt	<=	99	;
						10'd737	:	dt	<=	83	;
						10'd738	:	dt	<=	101	;
						10'd739	:	dt	<=	94	;
						10'd740	:	dt	<=	71	;
						10'd741	:	dt	<=	32	;
						10'd742	:	dt	<=	2	;
						10'd743	:	dt	<=	15	;
						10'd744	:	dt	<=	36	;
						10'd745	:	dt	<=	0	;
						10'd746	:	dt	<=	4	;
						10'd747	:	dt	<=	31	;
						10'd748	:	dt	<=	27	;
						10'd749	:	dt	<=	22	;
						10'd750	:	dt	<=	19	;
						10'd751	:	dt	<=	16	;
						10'd752	:	dt	<=	9	;
						10'd753	:	dt	<=	13	;
						10'd754	:	dt	<=	16	;
						10'd755	:	dt	<=	5	;
						10'd756	:	dt	<=	89	;
						10'd757	:	dt	<=	90	;
						10'd758	:	dt	<=	90	;
						10'd759	:	dt	<=	94	;
						10'd760	:	dt	<=	163	;
						10'd761	:	dt	<=	154	;
						10'd762	:	dt	<=	126	;
						10'd763	:	dt	<=	110	;
						10'd764	:	dt	<=	96	;
						10'd765	:	dt	<=	86	;
						10'd766	:	dt	<=	91	;
						10'd767	:	dt	<=	82	;
						10'd768	:	dt	<=	29	;
						10'd769	:	dt	<=	16	;
						10'd770	:	dt	<=	13	;
						10'd771	:	dt	<=	8	;
						10'd772	:	dt	<=	35	;
						10'd773	:	dt	<=	16	;
						10'd774	:	dt	<=	0	;
						10'd775	:	dt	<=	20	;
						10'd776	:	dt	<=	30	;
						10'd777	:	dt	<=	20	;
						10'd778	:	dt	<=	19	;
						10'd779	:	dt	<=	17	;
						10'd780	:	dt	<=	13	;
						10'd781	:	dt	<=	10	;
						10'd782	:	dt	<=	7	;
						10'd783	:	dt	<=	9	;
					endcase
				end
				5'd12	:	begin
					case (cnt)
						10'd0	:	dt	<=	178	;
						10'd1	:	dt	<=	179	;
						10'd2	:	dt	<=	181	;
						10'd3	:	dt	<=	183	;
						10'd4	:	dt	<=	184	;
						10'd5	:	dt	<=	183	;
						10'd6	:	dt	<=	183	;
						10'd7	:	dt	<=	184	;
						10'd8	:	dt	<=	185	;
						10'd9	:	dt	<=	186	;
						10'd10	:	dt	<=	185	;
						10'd11	:	dt	<=	184	;
						10'd12	:	dt	<=	184	;
						10'd13	:	dt	<=	183	;
						10'd14	:	dt	<=	185	;
						10'd15	:	dt	<=	187	;
						10'd16	:	dt	<=	182	;
						10'd17	:	dt	<=	179	;
						10'd18	:	dt	<=	179	;
						10'd19	:	dt	<=	177	;
						10'd20	:	dt	<=	177	;
						10'd21	:	dt	<=	177	;
						10'd22	:	dt	<=	174	;
						10'd23	:	dt	<=	173	;
						10'd24	:	dt	<=	172	;
						10'd25	:	dt	<=	170	;
						10'd26	:	dt	<=	169	;
						10'd27	:	dt	<=	166	;
						10'd28	:	dt	<=	179	;
						10'd29	:	dt	<=	184	;
						10'd30	:	dt	<=	185	;
						10'd31	:	dt	<=	185	;
						10'd32	:	dt	<=	186	;
						10'd33	:	dt	<=	187	;
						10'd34	:	dt	<=	186	;
						10'd35	:	dt	<=	186	;
						10'd36	:	dt	<=	187	;
						10'd37	:	dt	<=	187	;
						10'd38	:	dt	<=	188	;
						10'd39	:	dt	<=	188	;
						10'd40	:	dt	<=	186	;
						10'd41	:	dt	<=	185	;
						10'd42	:	dt	<=	174	;
						10'd43	:	dt	<=	158	;
						10'd44	:	dt	<=	171	;
						10'd45	:	dt	<=	185	;
						10'd46	:	dt	<=	179	;
						10'd47	:	dt	<=	179	;
						10'd48	:	dt	<=	179	;
						10'd49	:	dt	<=	177	;
						10'd50	:	dt	<=	175	;
						10'd51	:	dt	<=	174	;
						10'd52	:	dt	<=	174	;
						10'd53	:	dt	<=	172	;
						10'd54	:	dt	<=	169	;
						10'd55	:	dt	<=	167	;
						10'd56	:	dt	<=	182	;
						10'd57	:	dt	<=	184	;
						10'd58	:	dt	<=	185	;
						10'd59	:	dt	<=	187	;
						10'd60	:	dt	<=	187	;
						10'd61	:	dt	<=	188	;
						10'd62	:	dt	<=	189	;
						10'd63	:	dt	<=	189	;
						10'd64	:	dt	<=	188	;
						10'd65	:	dt	<=	188	;
						10'd66	:	dt	<=	187	;
						10'd67	:	dt	<=	173	;
						10'd68	:	dt	<=	184	;
						10'd69	:	dt	<=	188	;
						10'd70	:	dt	<=	135	;
						10'd71	:	dt	<=	105	;
						10'd72	:	dt	<=	82	;
						10'd73	:	dt	<=	160	;
						10'd74	:	dt	<=	191	;
						10'd75	:	dt	<=	183	;
						10'd76	:	dt	<=	184	;
						10'd77	:	dt	<=	181	;
						10'd78	:	dt	<=	176	;
						10'd79	:	dt	<=	176	;
						10'd80	:	dt	<=	175	;
						10'd81	:	dt	<=	175	;
						10'd82	:	dt	<=	171	;
						10'd83	:	dt	<=	169	;
						10'd84	:	dt	<=	184	;
						10'd85	:	dt	<=	186	;
						10'd86	:	dt	<=	187	;
						10'd87	:	dt	<=	188	;
						10'd88	:	dt	<=	188	;
						10'd89	:	dt	<=	188	;
						10'd90	:	dt	<=	189	;
						10'd91	:	dt	<=	191	;
						10'd92	:	dt	<=	188	;
						10'd93	:	dt	<=	190	;
						10'd94	:	dt	<=	169	;
						10'd95	:	dt	<=	118	;
						10'd96	:	dt	<=	98	;
						10'd97	:	dt	<=	145	;
						10'd98	:	dt	<=	147	;
						10'd99	:	dt	<=	120	;
						10'd100	:	dt	<=	80	;
						10'd101	:	dt	<=	89	;
						10'd102	:	dt	<=	170	;
						10'd103	:	dt	<=	132	;
						10'd104	:	dt	<=	118	;
						10'd105	:	dt	<=	157	;
						10'd106	:	dt	<=	184	;
						10'd107	:	dt	<=	175	;
						10'd108	:	dt	<=	175	;
						10'd109	:	dt	<=	174	;
						10'd110	:	dt	<=	172	;
						10'd111	:	dt	<=	170	;
						10'd112	:	dt	<=	186	;
						10'd113	:	dt	<=	188	;
						10'd114	:	dt	<=	188	;
						10'd115	:	dt	<=	188	;
						10'd116	:	dt	<=	189	;
						10'd117	:	dt	<=	192	;
						10'd118	:	dt	<=	190	;
						10'd119	:	dt	<=	190	;
						10'd120	:	dt	<=	188	;
						10'd121	:	dt	<=	199	;
						10'd122	:	dt	<=	167	;
						10'd123	:	dt	<=	133	;
						10'd124	:	dt	<=	93	;
						10'd125	:	dt	<=	83	;
						10'd126	:	dt	<=	164	;
						10'd127	:	dt	<=	129	;
						10'd128	:	dt	<=	103	;
						10'd129	:	dt	<=	76	;
						10'd130	:	dt	<=	74	;
						10'd131	:	dt	<=	104	;
						10'd132	:	dt	<=	86	;
						10'd133	:	dt	<=	61	;
						10'd134	:	dt	<=	157	;
						10'd135	:	dt	<=	185	;
						10'd136	:	dt	<=	177	;
						10'd137	:	dt	<=	175	;
						10'd138	:	dt	<=	173	;
						10'd139	:	dt	<=	171	;
						10'd140	:	dt	<=	186	;
						10'd141	:	dt	<=	187	;
						10'd142	:	dt	<=	189	;
						10'd143	:	dt	<=	189	;
						10'd144	:	dt	<=	191	;
						10'd145	:	dt	<=	191	;
						10'd146	:	dt	<=	193	;
						10'd147	:	dt	<=	193	;
						10'd148	:	dt	<=	190	;
						10'd149	:	dt	<=	203	;
						10'd150	:	dt	<=	179	;
						10'd151	:	dt	<=	148	;
						10'd152	:	dt	<=	124	;
						10'd153	:	dt	<=	73	;
						10'd154	:	dt	<=	158	;
						10'd155	:	dt	<=	142	;
						10'd156	:	dt	<=	111	;
						10'd157	:	dt	<=	83	;
						10'd158	:	dt	<=	51	;
						10'd159	:	dt	<=	98	;
						10'd160	:	dt	<=	94	;
						10'd161	:	dt	<=	42	;
						10'd162	:	dt	<=	87	;
						10'd163	:	dt	<=	192	;
						10'd164	:	dt	<=	178	;
						10'd165	:	dt	<=	177	;
						10'd166	:	dt	<=	175	;
						10'd167	:	dt	<=	172	;
						10'd168	:	dt	<=	187	;
						10'd169	:	dt	<=	189	;
						10'd170	:	dt	<=	189	;
						10'd171	:	dt	<=	190	;
						10'd172	:	dt	<=	192	;
						10'd173	:	dt	<=	192	;
						10'd174	:	dt	<=	193	;
						10'd175	:	dt	<=	192	;
						10'd176	:	dt	<=	197	;
						10'd177	:	dt	<=	206	;
						10'd178	:	dt	<=	196	;
						10'd179	:	dt	<=	157	;
						10'd180	:	dt	<=	130	;
						10'd181	:	dt	<=	76	;
						10'd182	:	dt	<=	127	;
						10'd183	:	dt	<=	148	;
						10'd184	:	dt	<=	114	;
						10'd185	:	dt	<=	88	;
						10'd186	:	dt	<=	40	;
						10'd187	:	dt	<=	93	;
						10'd188	:	dt	<=	90	;
						10'd189	:	dt	<=	51	;
						10'd190	:	dt	<=	57	;
						10'd191	:	dt	<=	189	;
						10'd192	:	dt	<=	179	;
						10'd193	:	dt	<=	178	;
						10'd194	:	dt	<=	177	;
						10'd195	:	dt	<=	175	;
						10'd196	:	dt	<=	190	;
						10'd197	:	dt	<=	192	;
						10'd198	:	dt	<=	191	;
						10'd199	:	dt	<=	192	;
						10'd200	:	dt	<=	193	;
						10'd201	:	dt	<=	193	;
						10'd202	:	dt	<=	194	;
						10'd203	:	dt	<=	192	;
						10'd204	:	dt	<=	205	;
						10'd205	:	dt	<=	182	;
						10'd206	:	dt	<=	205	;
						10'd207	:	dt	<=	165	;
						10'd208	:	dt	<=	132	;
						10'd209	:	dt	<=	85	;
						10'd210	:	dt	<=	93	;
						10'd211	:	dt	<=	148	;
						10'd212	:	dt	<=	116	;
						10'd213	:	dt	<=	89	;
						10'd214	:	dt	<=	41	;
						10'd215	:	dt	<=	78	;
						10'd216	:	dt	<=	98	;
						10'd217	:	dt	<=	53	;
						10'd218	:	dt	<=	60	;
						10'd219	:	dt	<=	190	;
						10'd220	:	dt	<=	179	;
						10'd221	:	dt	<=	179	;
						10'd222	:	dt	<=	177	;
						10'd223	:	dt	<=	176	;
						10'd224	:	dt	<=	190	;
						10'd225	:	dt	<=	191	;
						10'd226	:	dt	<=	192	;
						10'd227	:	dt	<=	192	;
						10'd228	:	dt	<=	192	;
						10'd229	:	dt	<=	194	;
						10'd230	:	dt	<=	191	;
						10'd231	:	dt	<=	189	;
						10'd232	:	dt	<=	178	;
						10'd233	:	dt	<=	113	;
						10'd234	:	dt	<=	164	;
						10'd235	:	dt	<=	174	;
						10'd236	:	dt	<=	123	;
						10'd237	:	dt	<=	93	;
						10'd238	:	dt	<=	77	;
						10'd239	:	dt	<=	149	;
						10'd240	:	dt	<=	119	;
						10'd241	:	dt	<=	93	;
						10'd242	:	dt	<=	49	;
						10'd243	:	dt	<=	68	;
						10'd244	:	dt	<=	101	;
						10'd245	:	dt	<=	51	;
						10'd246	:	dt	<=	78	;
						10'd247	:	dt	<=	195	;
						10'd248	:	dt	<=	179	;
						10'd249	:	dt	<=	181	;
						10'd250	:	dt	<=	179	;
						10'd251	:	dt	<=	178	;
						10'd252	:	dt	<=	189	;
						10'd253	:	dt	<=	191	;
						10'd254	:	dt	<=	192	;
						10'd255	:	dt	<=	193	;
						10'd256	:	dt	<=	194	;
						10'd257	:	dt	<=	190	;
						10'd258	:	dt	<=	189	;
						10'd259	:	dt	<=	196	;
						10'd260	:	dt	<=	159	;
						10'd261	:	dt	<=	93	;
						10'd262	:	dt	<=	83	;
						10'd263	:	dt	<=	167	;
						10'd264	:	dt	<=	129	;
						10'd265	:	dt	<=	92	;
						10'd266	:	dt	<=	55	;
						10'd267	:	dt	<=	143	;
						10'd268	:	dt	<=	133	;
						10'd269	:	dt	<=	100	;
						10'd270	:	dt	<=	63	;
						10'd271	:	dt	<=	42	;
						10'd272	:	dt	<=	83	;
						10'd273	:	dt	<=	43	;
						10'd274	:	dt	<=	121	;
						10'd275	:	dt	<=	197	;
						10'd276	:	dt	<=	181	;
						10'd277	:	dt	<=	182	;
						10'd278	:	dt	<=	181	;
						10'd279	:	dt	<=	179	;
						10'd280	:	dt	<=	191	;
						10'd281	:	dt	<=	193	;
						10'd282	:	dt	<=	194	;
						10'd283	:	dt	<=	194	;
						10'd284	:	dt	<=	194	;
						10'd285	:	dt	<=	206	;
						10'd286	:	dt	<=	206	;
						10'd287	:	dt	<=	182	;
						10'd288	:	dt	<=	130	;
						10'd289	:	dt	<=	91	;
						10'd290	:	dt	<=	51	;
						10'd291	:	dt	<=	138	;
						10'd292	:	dt	<=	133	;
						10'd293	:	dt	<=	80	;
						10'd294	:	dt	<=	43	;
						10'd295	:	dt	<=	131	;
						10'd296	:	dt	<=	165	;
						10'd297	:	dt	<=	126	;
						10'd298	:	dt	<=	79	;
						10'd299	:	dt	<=	38	;
						10'd300	:	dt	<=	64	;
						10'd301	:	dt	<=	35	;
						10'd302	:	dt	<=	143	;
						10'd303	:	dt	<=	195	;
						10'd304	:	dt	<=	183	;
						10'd305	:	dt	<=	184	;
						10'd306	:	dt	<=	181	;
						10'd307	:	dt	<=	179	;
						10'd308	:	dt	<=	192	;
						10'd309	:	dt	<=	193	;
						10'd310	:	dt	<=	196	;
						10'd311	:	dt	<=	194	;
						10'd312	:	dt	<=	203	;
						10'd313	:	dt	<=	204	;
						10'd314	:	dt	<=	177	;
						10'd315	:	dt	<=	163	;
						10'd316	:	dt	<=	119	;
						10'd317	:	dt	<=	105	;
						10'd318	:	dt	<=	56	;
						10'd319	:	dt	<=	112	;
						10'd320	:	dt	<=	134	;
						10'd321	:	dt	<=	92	;
						10'd322	:	dt	<=	56	;
						10'd323	:	dt	<=	141	;
						10'd324	:	dt	<=	183	;
						10'd325	:	dt	<=	134	;
						10'd326	:	dt	<=	82	;
						10'd327	:	dt	<=	48	;
						10'd328	:	dt	<=	73	;
						10'd329	:	dt	<=	53	;
						10'd330	:	dt	<=	168	;
						10'd331	:	dt	<=	192	;
						10'd332	:	dt	<=	186	;
						10'd333	:	dt	<=	184	;
						10'd334	:	dt	<=	182	;
						10'd335	:	dt	<=	181	;
						10'd336	:	dt	<=	193	;
						10'd337	:	dt	<=	194	;
						10'd338	:	dt	<=	195	;
						10'd339	:	dt	<=	194	;
						10'd340	:	dt	<=	218	;
						10'd341	:	dt	<=	193	;
						10'd342	:	dt	<=	145	;
						10'd343	:	dt	<=	164	;
						10'd344	:	dt	<=	128	;
						10'd345	:	dt	<=	115	;
						10'd346	:	dt	<=	66	;
						10'd347	:	dt	<=	78	;
						10'd348	:	dt	<=	147	;
						10'd349	:	dt	<=	133	;
						10'd350	:	dt	<=	78	;
						10'd351	:	dt	<=	105	;
						10'd352	:	dt	<=	159	;
						10'd353	:	dt	<=	107	;
						10'd354	:	dt	<=	57	;
						10'd355	:	dt	<=	47	;
						10'd356	:	dt	<=	80	;
						10'd357	:	dt	<=	49	;
						10'd358	:	dt	<=	150	;
						10'd359	:	dt	<=	199	;
						10'd360	:	dt	<=	186	;
						10'd361	:	dt	<=	184	;
						10'd362	:	dt	<=	183	;
						10'd363	:	dt	<=	180	;
						10'd364	:	dt	<=	194	;
						10'd365	:	dt	<=	194	;
						10'd366	:	dt	<=	193	;
						10'd367	:	dt	<=	203	;
						10'd368	:	dt	<=	199	;
						10'd369	:	dt	<=	171	;
						10'd370	:	dt	<=	124	;
						10'd371	:	dt	<=	122	;
						10'd372	:	dt	<=	139	;
						10'd373	:	dt	<=	108	;
						10'd374	:	dt	<=	67	;
						10'd375	:	dt	<=	52	;
						10'd376	:	dt	<=	154	;
						10'd377	:	dt	<=	144	;
						10'd378	:	dt	<=	106	;
						10'd379	:	dt	<=	38	;
						10'd380	:	dt	<=	36	;
						10'd381	:	dt	<=	35	;
						10'd382	:	dt	<=	30	;
						10'd383	:	dt	<=	69	;
						10'd384	:	dt	<=	79	;
						10'd385	:	dt	<=	28	;
						10'd386	:	dt	<=	75	;
						10'd387	:	dt	<=	202	;
						10'd388	:	dt	<=	186	;
						10'd389	:	dt	<=	186	;
						10'd390	:	dt	<=	185	;
						10'd391	:	dt	<=	182	;
						10'd392	:	dt	<=	195	;
						10'd393	:	dt	<=	195	;
						10'd394	:	dt	<=	195	;
						10'd395	:	dt	<=	204	;
						10'd396	:	dt	<=	188	;
						10'd397	:	dt	<=	154	;
						10'd398	:	dt	<=	125	;
						10'd399	:	dt	<=	80	;
						10'd400	:	dt	<=	121	;
						10'd401	:	dt	<=	116	;
						10'd402	:	dt	<=	88	;
						10'd403	:	dt	<=	42	;
						10'd404	:	dt	<=	126	;
						10'd405	:	dt	<=	144	;
						10'd406	:	dt	<=	96	;
						10'd407	:	dt	<=	41	;
						10'd408	:	dt	<=	16	;
						10'd409	:	dt	<=	55	;
						10'd410	:	dt	<=	67	;
						10'd411	:	dt	<=	67	;
						10'd412	:	dt	<=	46	;
						10'd413	:	dt	<=	38	;
						10'd414	:	dt	<=	43	;
						10'd415	:	dt	<=	184	;
						10'd416	:	dt	<=	192	;
						10'd417	:	dt	<=	187	;
						10'd418	:	dt	<=	185	;
						10'd419	:	dt	<=	183	;
						10'd420	:	dt	<=	192	;
						10'd421	:	dt	<=	196	;
						10'd422	:	dt	<=	197	;
						10'd423	:	dt	<=	200	;
						10'd424	:	dt	<=	202	;
						10'd425	:	dt	<=	173	;
						10'd426	:	dt	<=	144	;
						10'd427	:	dt	<=	103	;
						10'd428	:	dt	<=	86	;
						10'd429	:	dt	<=	130	;
						10'd430	:	dt	<=	89	;
						10'd431	:	dt	<=	48	;
						10'd432	:	dt	<=	25	;
						10'd433	:	dt	<=	85	;
						10'd434	:	dt	<=	89	;
						10'd435	:	dt	<=	44	;
						10'd436	:	dt	<=	70	;
						10'd437	:	dt	<=	97	;
						10'd438	:	dt	<=	113	;
						10'd439	:	dt	<=	92	;
						10'd440	:	dt	<=	58	;
						10'd441	:	dt	<=	45	;
						10'd442	:	dt	<=	59	;
						10'd443	:	dt	<=	190	;
						10'd444	:	dt	<=	189	;
						10'd445	:	dt	<=	188	;
						10'd446	:	dt	<=	185	;
						10'd447	:	dt	<=	185	;
						10'd448	:	dt	<=	194	;
						10'd449	:	dt	<=	197	;
						10'd450	:	dt	<=	198	;
						10'd451	:	dt	<=	201	;
						10'd452	:	dt	<=	206	;
						10'd453	:	dt	<=	180	;
						10'd454	:	dt	<=	149	;
						10'd455	:	dt	<=	119	;
						10'd456	:	dt	<=	81	;
						10'd457	:	dt	<=	106	;
						10'd458	:	dt	<=	81	;
						10'd459	:	dt	<=	70	;
						10'd460	:	dt	<=	20	;
						10'd461	:	dt	<=	92	;
						10'd462	:	dt	<=	164	;
						10'd463	:	dt	<=	137	;
						10'd464	:	dt	<=	127	;
						10'd465	:	dt	<=	116	;
						10'd466	:	dt	<=	124	;
						10'd467	:	dt	<=	98	;
						10'd468	:	dt	<=	66	;
						10'd469	:	dt	<=	26	;
						10'd470	:	dt	<=	111	;
						10'd471	:	dt	<=	205	;
						10'd472	:	dt	<=	188	;
						10'd473	:	dt	<=	190	;
						10'd474	:	dt	<=	186	;
						10'd475	:	dt	<=	184	;
						10'd476	:	dt	<=	196	;
						10'd477	:	dt	<=	197	;
						10'd478	:	dt	<=	200	;
						10'd479	:	dt	<=	202	;
						10'd480	:	dt	<=	208	;
						10'd481	:	dt	<=	190	;
						10'd482	:	dt	<=	158	;
						10'd483	:	dt	<=	130	;
						10'd484	:	dt	<=	98	;
						10'd485	:	dt	<=	74	;
						10'd486	:	dt	<=	95	;
						10'd487	:	dt	<=	103	;
						10'd488	:	dt	<=	63	;
						10'd489	:	dt	<=	158	;
						10'd490	:	dt	<=	196	;
						10'd491	:	dt	<=	177	;
						10'd492	:	dt	<=	148	;
						10'd493	:	dt	<=	125	;
						10'd494	:	dt	<=	117	;
						10'd495	:	dt	<=	89	;
						10'd496	:	dt	<=	58	;
						10'd497	:	dt	<=	22	;
						10'd498	:	dt	<=	153	;
						10'd499	:	dt	<=	203	;
						10'd500	:	dt	<=	190	;
						10'd501	:	dt	<=	190	;
						10'd502	:	dt	<=	187	;
						10'd503	:	dt	<=	184	;
						10'd504	:	dt	<=	195	;
						10'd505	:	dt	<=	197	;
						10'd506	:	dt	<=	199	;
						10'd507	:	dt	<=	205	;
						10'd508	:	dt	<=	200	;
						10'd509	:	dt	<=	180	;
						10'd510	:	dt	<=	155	;
						10'd511	:	dt	<=	128	;
						10'd512	:	dt	<=	98	;
						10'd513	:	dt	<=	76	;
						10'd514	:	dt	<=	83	;
						10'd515	:	dt	<=	99	;
						10'd516	:	dt	<=	121	;
						10'd517	:	dt	<=	191	;
						10'd518	:	dt	<=	186	;
						10'd519	:	dt	<=	165	;
						10'd520	:	dt	<=	140	;
						10'd521	:	dt	<=	121	;
						10'd522	:	dt	<=	102	;
						10'd523	:	dt	<=	84	;
						10'd524	:	dt	<=	47	;
						10'd525	:	dt	<=	31	;
						10'd526	:	dt	<=	182	;
						10'd527	:	dt	<=	196	;
						10'd528	:	dt	<=	192	;
						10'd529	:	dt	<=	190	;
						10'd530	:	dt	<=	187	;
						10'd531	:	dt	<=	186	;
						10'd532	:	dt	<=	197	;
						10'd533	:	dt	<=	199	;
						10'd534	:	dt	<=	201	;
						10'd535	:	dt	<=	202	;
						10'd536	:	dt	<=	186	;
						10'd537	:	dt	<=	169	;
						10'd538	:	dt	<=	155	;
						10'd539	:	dt	<=	128	;
						10'd540	:	dt	<=	91	;
						10'd541	:	dt	<=	103	;
						10'd542	:	dt	<=	73	;
						10'd543	:	dt	<=	109	;
						10'd544	:	dt	<=	173	;
						10'd545	:	dt	<=	183	;
						10'd546	:	dt	<=	174	;
						10'd547	:	dt	<=	153	;
						10'd548	:	dt	<=	132	;
						10'd549	:	dt	<=	114	;
						10'd550	:	dt	<=	94	;
						10'd551	:	dt	<=	79	;
						10'd552	:	dt	<=	29	;
						10'd553	:	dt	<=	91	;
						10'd554	:	dt	<=	207	;
						10'd555	:	dt	<=	190	;
						10'd556	:	dt	<=	192	;
						10'd557	:	dt	<=	190	;
						10'd558	:	dt	<=	188	;
						10'd559	:	dt	<=	187	;
						10'd560	:	dt	<=	197	;
						10'd561	:	dt	<=	200	;
						10'd562	:	dt	<=	201	;
						10'd563	:	dt	<=	199	;
						10'd564	:	dt	<=	186	;
						10'd565	:	dt	<=	173	;
						10'd566	:	dt	<=	159	;
						10'd567	:	dt	<=	124	;
						10'd568	:	dt	<=	94	;
						10'd569	:	dt	<=	117	;
						10'd570	:	dt	<=	97	;
						10'd571	:	dt	<=	159	;
						10'd572	:	dt	<=	177	;
						10'd573	:	dt	<=	175	;
						10'd574	:	dt	<=	167	;
						10'd575	:	dt	<=	143	;
						10'd576	:	dt	<=	123	;
						10'd577	:	dt	<=	103	;
						10'd578	:	dt	<=	85	;
						10'd579	:	dt	<=	55	;
						10'd580	:	dt	<=	45	;
						10'd581	:	dt	<=	187	;
						10'd582	:	dt	<=	198	;
						10'd583	:	dt	<=	193	;
						10'd584	:	dt	<=	192	;
						10'd585	:	dt	<=	191	;
						10'd586	:	dt	<=	188	;
						10'd587	:	dt	<=	187	;
						10'd588	:	dt	<=	199	;
						10'd589	:	dt	<=	201	;
						10'd590	:	dt	<=	201	;
						10'd591	:	dt	<=	203	;
						10'd592	:	dt	<=	190	;
						10'd593	:	dt	<=	171	;
						10'd594	:	dt	<=	160	;
						10'd595	:	dt	<=	131	;
						10'd596	:	dt	<=	110	;
						10'd597	:	dt	<=	107	;
						10'd598	:	dt	<=	109	;
						10'd599	:	dt	<=	166	;
						10'd600	:	dt	<=	165	;
						10'd601	:	dt	<=	173	;
						10'd602	:	dt	<=	162	;
						10'd603	:	dt	<=	136	;
						10'd604	:	dt	<=	109	;
						10'd605	:	dt	<=	89	;
						10'd606	:	dt	<=	78	;
						10'd607	:	dt	<=	29	;
						10'd608	:	dt	<=	103	;
						10'd609	:	dt	<=	214	;
						10'd610	:	dt	<=	194	;
						10'd611	:	dt	<=	195	;
						10'd612	:	dt	<=	193	;
						10'd613	:	dt	<=	193	;
						10'd614	:	dt	<=	191	;
						10'd615	:	dt	<=	188	;
						10'd616	:	dt	<=	198	;
						10'd617	:	dt	<=	201	;
						10'd618	:	dt	<=	201	;
						10'd619	:	dt	<=	204	;
						10'd620	:	dt	<=	193	;
						10'd621	:	dt	<=	175	;
						10'd622	:	dt	<=	163	;
						10'd623	:	dt	<=	142	;
						10'd624	:	dt	<=	118	;
						10'd625	:	dt	<=	93	;
						10'd626	:	dt	<=	107	;
						10'd627	:	dt	<=	163	;
						10'd628	:	dt	<=	159	;
						10'd629	:	dt	<=	162	;
						10'd630	:	dt	<=	145	;
						10'd631	:	dt	<=	123	;
						10'd632	:	dt	<=	94	;
						10'd633	:	dt	<=	77	;
						10'd634	:	dt	<=	59	;
						10'd635	:	dt	<=	23	;
						10'd636	:	dt	<=	174	;
						10'd637	:	dt	<=	206	;
						10'd638	:	dt	<=	199	;
						10'd639	:	dt	<=	196	;
						10'd640	:	dt	<=	194	;
						10'd641	:	dt	<=	193	;
						10'd642	:	dt	<=	192	;
						10'd643	:	dt	<=	190	;
						10'd644	:	dt	<=	198	;
						10'd645	:	dt	<=	201	;
						10'd646	:	dt	<=	202	;
						10'd647	:	dt	<=	203	;
						10'd648	:	dt	<=	200	;
						10'd649	:	dt	<=	187	;
						10'd650	:	dt	<=	164	;
						10'd651	:	dt	<=	139	;
						10'd652	:	dt	<=	116	;
						10'd653	:	dt	<=	88	;
						10'd654	:	dt	<=	98	;
						10'd655	:	dt	<=	148	;
						10'd656	:	dt	<=	148	;
						10'd657	:	dt	<=	142	;
						10'd658	:	dt	<=	127	;
						10'd659	:	dt	<=	101	;
						10'd660	:	dt	<=	77	;
						10'd661	:	dt	<=	67	;
						10'd662	:	dt	<=	26	;
						10'd663	:	dt	<=	84	;
						10'd664	:	dt	<=	214	;
						10'd665	:	dt	<=	200	;
						10'd666	:	dt	<=	198	;
						10'd667	:	dt	<=	196	;
						10'd668	:	dt	<=	194	;
						10'd669	:	dt	<=	193	;
						10'd670	:	dt	<=	192	;
						10'd671	:	dt	<=	191	;
						10'd672	:	dt	<=	198	;
						10'd673	:	dt	<=	201	;
						10'd674	:	dt	<=	203	;
						10'd675	:	dt	<=	203	;
						10'd676	:	dt	<=	203	;
						10'd677	:	dt	<=	185	;
						10'd678	:	dt	<=	161	;
						10'd679	:	dt	<=	142	;
						10'd680	:	dt	<=	121	;
						10'd681	:	dt	<=	102	;
						10'd682	:	dt	<=	100	;
						10'd683	:	dt	<=	134	;
						10'd684	:	dt	<=	137	;
						10'd685	:	dt	<=	120	;
						10'd686	:	dt	<=	106	;
						10'd687	:	dt	<=	88	;
						10'd688	:	dt	<=	68	;
						10'd689	:	dt	<=	45	;
						10'd690	:	dt	<=	30	;
						10'd691	:	dt	<=	185	;
						10'd692	:	dt	<=	206	;
						10'd693	:	dt	<=	199	;
						10'd694	:	dt	<=	198	;
						10'd695	:	dt	<=	195	;
						10'd696	:	dt	<=	195	;
						10'd697	:	dt	<=	194	;
						10'd698	:	dt	<=	193	;
						10'd699	:	dt	<=	191	;
						10'd700	:	dt	<=	200	;
						10'd701	:	dt	<=	201	;
						10'd702	:	dt	<=	204	;
						10'd703	:	dt	<=	203	;
						10'd704	:	dt	<=	206	;
						10'd705	:	dt	<=	177	;
						10'd706	:	dt	<=	148	;
						10'd707	:	dt	<=	134	;
						10'd708	:	dt	<=	116	;
						10'd709	:	dt	<=	113	;
						10'd710	:	dt	<=	103	;
						10'd711	:	dt	<=	124	;
						10'd712	:	dt	<=	140	;
						10'd713	:	dt	<=	121	;
						10'd714	:	dt	<=	101	;
						10'd715	:	dt	<=	83	;
						10'd716	:	dt	<=	64	;
						10'd717	:	dt	<=	16	;
						10'd718	:	dt	<=	132	;
						10'd719	:	dt	<=	215	;
						10'd720	:	dt	<=	199	;
						10'd721	:	dt	<=	200	;
						10'd722	:	dt	<=	199	;
						10'd723	:	dt	<=	197	;
						10'd724	:	dt	<=	194	;
						10'd725	:	dt	<=	194	;
						10'd726	:	dt	<=	195	;
						10'd727	:	dt	<=	192	;
						10'd728	:	dt	<=	201	;
						10'd729	:	dt	<=	202	;
						10'd730	:	dt	<=	204	;
						10'd731	:	dt	<=	203	;
						10'd732	:	dt	<=	206	;
						10'd733	:	dt	<=	175	;
						10'd734	:	dt	<=	151	;
						10'd735	:	dt	<=	142	;
						10'd736	:	dt	<=	134	;
						10'd737	:	dt	<=	132	;
						10'd738	:	dt	<=	118	;
						10'd739	:	dt	<=	124	;
						10'd740	:	dt	<=	136	;
						10'd741	:	dt	<=	118	;
						10'd742	:	dt	<=	96	;
						10'd743	:	dt	<=	76	;
						10'd744	:	dt	<=	38	;
						10'd745	:	dt	<=	68	;
						10'd746	:	dt	<=	211	;
						10'd747	:	dt	<=	203	;
						10'd748	:	dt	<=	203	;
						10'd749	:	dt	<=	201	;
						10'd750	:	dt	<=	199	;
						10'd751	:	dt	<=	199	;
						10'd752	:	dt	<=	196	;
						10'd753	:	dt	<=	194	;
						10'd754	:	dt	<=	194	;
						10'd755	:	dt	<=	193	;
						10'd756	:	dt	<=	201	;
						10'd757	:	dt	<=	202	;
						10'd758	:	dt	<=	203	;
						10'd759	:	dt	<=	198	;
						10'd760	:	dt	<=	202	;
						10'd761	:	dt	<=	177	;
						10'd762	:	dt	<=	156	;
						10'd763	:	dt	<=	156	;
						10'd764	:	dt	<=	147	;
						10'd765	:	dt	<=	135	;
						10'd766	:	dt	<=	125	;
						10'd767	:	dt	<=	126	;
						10'd768	:	dt	<=	132	;
						10'd769	:	dt	<=	111	;
						10'd770	:	dt	<=	73	;
						10'd771	:	dt	<=	61	;
						10'd772	:	dt	<=	29	;
						10'd773	:	dt	<=	156	;
						10'd774	:	dt	<=	215	;
						10'd775	:	dt	<=	202	;
						10'd776	:	dt	<=	204	;
						10'd777	:	dt	<=	202	;
						10'd778	:	dt	<=	201	;
						10'd779	:	dt	<=	200	;
						10'd780	:	dt	<=	198	;
						10'd781	:	dt	<=	196	;
						10'd782	:	dt	<=	194	;
						10'd783	:	dt	<=	193	;
					endcase
				end
				5'd13	:	begin
					case (cnt)	
						10'd0	:	dt	<=	167	;
						10'd1	:	dt	<=	169	;
						10'd2	:	dt	<=	173	;
						10'd3	:	dt	<=	180	;
						10'd4	:	dt	<=	186	;
						10'd5	:	dt	<=	189	;
						10'd6	:	dt	<=	192	;
						10'd7	:	dt	<=	193	;
						10'd8	:	dt	<=	196	;
						10'd9	:	dt	<=	199	;
						10'd10	:	dt	<=	203	;
						10'd11	:	dt	<=	205	;
						10'd12	:	dt	<=	206	;
						10'd13	:	dt	<=	208	;
						10'd14	:	dt	<=	210	;
						10'd15	:	dt	<=	211	;
						10'd16	:	dt	<=	212	;
						10'd17	:	dt	<=	213	;
						10'd18	:	dt	<=	212	;
						10'd19	:	dt	<=	214	;
						10'd20	:	dt	<=	215	;
						10'd21	:	dt	<=	213	;
						10'd22	:	dt	<=	214	;
						10'd23	:	dt	<=	213	;
						10'd24	:	dt	<=	214	;
						10'd25	:	dt	<=	215	;
						10'd26	:	dt	<=	214	;
						10'd27	:	dt	<=	213	;
						10'd28	:	dt	<=	169	;
						10'd29	:	dt	<=	171	;
						10'd30	:	dt	<=	175	;
						10'd31	:	dt	<=	181	;
						10'd32	:	dt	<=	187	;
						10'd33	:	dt	<=	190	;
						10'd34	:	dt	<=	193	;
						10'd35	:	dt	<=	194	;
						10'd36	:	dt	<=	197	;
						10'd37	:	dt	<=	200	;
						10'd38	:	dt	<=	203	;
						10'd39	:	dt	<=	206	;
						10'd40	:	dt	<=	207	;
						10'd41	:	dt	<=	210	;
						10'd42	:	dt	<=	212	;
						10'd43	:	dt	<=	212	;
						10'd44	:	dt	<=	213	;
						10'd45	:	dt	<=	214	;
						10'd46	:	dt	<=	214	;
						10'd47	:	dt	<=	216	;
						10'd48	:	dt	<=	216	;
						10'd49	:	dt	<=	215	;
						10'd50	:	dt	<=	215	;
						10'd51	:	dt	<=	215	;
						10'd52	:	dt	<=	217	;
						10'd53	:	dt	<=	217	;
						10'd54	:	dt	<=	217	;
						10'd55	:	dt	<=	215	;
						10'd56	:	dt	<=	171	;
						10'd57	:	dt	<=	173	;
						10'd58	:	dt	<=	177	;
						10'd59	:	dt	<=	183	;
						10'd60	:	dt	<=	190	;
						10'd61	:	dt	<=	192	;
						10'd62	:	dt	<=	194	;
						10'd63	:	dt	<=	196	;
						10'd64	:	dt	<=	199	;
						10'd65	:	dt	<=	202	;
						10'd66	:	dt	<=	204	;
						10'd67	:	dt	<=	207	;
						10'd68	:	dt	<=	209	;
						10'd69	:	dt	<=	212	;
						10'd70	:	dt	<=	213	;
						10'd71	:	dt	<=	214	;
						10'd72	:	dt	<=	214	;
						10'd73	:	dt	<=	216	;
						10'd74	:	dt	<=	216	;
						10'd75	:	dt	<=	215	;
						10'd76	:	dt	<=	216	;
						10'd77	:	dt	<=	216	;
						10'd78	:	dt	<=	218	;
						10'd79	:	dt	<=	217	;
						10'd80	:	dt	<=	218	;
						10'd81	:	dt	<=	218	;
						10'd82	:	dt	<=	218	;
						10'd83	:	dt	<=	217	;
						10'd84	:	dt	<=	173	;
						10'd85	:	dt	<=	175	;
						10'd86	:	dt	<=	180	;
						10'd87	:	dt	<=	185	;
						10'd88	:	dt	<=	191	;
						10'd89	:	dt	<=	194	;
						10'd90	:	dt	<=	197	;
						10'd91	:	dt	<=	199	;
						10'd92	:	dt	<=	201	;
						10'd93	:	dt	<=	204	;
						10'd94	:	dt	<=	206	;
						10'd95	:	dt	<=	208	;
						10'd96	:	dt	<=	211	;
						10'd97	:	dt	<=	213	;
						10'd98	:	dt	<=	214	;
						10'd99	:	dt	<=	212	;
						10'd100	:	dt	<=	215	;
						10'd101	:	dt	<=	211	;
						10'd102	:	dt	<=	215	;
						10'd103	:	dt	<=	223	;
						10'd104	:	dt	<=	223	;
						10'd105	:	dt	<=	220	;
						10'd106	:	dt	<=	218	;
						10'd107	:	dt	<=	219	;
						10'd108	:	dt	<=	220	;
						10'd109	:	dt	<=	219	;
						10'd110	:	dt	<=	218	;
						10'd111	:	dt	<=	218	;
						10'd112	:	dt	<=	175	;
						10'd113	:	dt	<=	176	;
						10'd114	:	dt	<=	181	;
						10'd115	:	dt	<=	187	;
						10'd116	:	dt	<=	191	;
						10'd117	:	dt	<=	195	;
						10'd118	:	dt	<=	198	;
						10'd119	:	dt	<=	201	;
						10'd120	:	dt	<=	204	;
						10'd121	:	dt	<=	206	;
						10'd122	:	dt	<=	208	;
						10'd123	:	dt	<=	210	;
						10'd124	:	dt	<=	213	;
						10'd125	:	dt	<=	214	;
						10'd126	:	dt	<=	220	;
						10'd127	:	dt	<=	240	;
						10'd128	:	dt	<=	238	;
						10'd129	:	dt	<=	200	;
						10'd130	:	dt	<=	162	;
						10'd131	:	dt	<=	196	;
						10'd132	:	dt	<=	209	;
						10'd133	:	dt	<=	219	;
						10'd134	:	dt	<=	225	;
						10'd135	:	dt	<=	220	;
						10'd136	:	dt	<=	221	;
						10'd137	:	dt	<=	221	;
						10'd138	:	dt	<=	220	;
						10'd139	:	dt	<=	220	;
						10'd140	:	dt	<=	176	;
						10'd141	:	dt	<=	178	;
						10'd142	:	dt	<=	183	;
						10'd143	:	dt	<=	189	;
						10'd144	:	dt	<=	193	;
						10'd145	:	dt	<=	197	;
						10'd146	:	dt	<=	200	;
						10'd147	:	dt	<=	203	;
						10'd148	:	dt	<=	205	;
						10'd149	:	dt	<=	207	;
						10'd150	:	dt	<=	211	;
						10'd151	:	dt	<=	211	;
						10'd152	:	dt	<=	214	;
						10'd153	:	dt	<=	213	;
						10'd154	:	dt	<=	214	;
						10'd155	:	dt	<=	232	;
						10'd156	:	dt	<=	242	;
						10'd157	:	dt	<=	199	;
						10'd158	:	dt	<=	145	;
						10'd159	:	dt	<=	123	;
						10'd160	:	dt	<=	163	;
						10'd161	:	dt	<=	165	;
						10'd162	:	dt	<=	201	;
						10'd163	:	dt	<=	226	;
						10'd164	:	dt	<=	221	;
						10'd165	:	dt	<=	222	;
						10'd166	:	dt	<=	222	;
						10'd167	:	dt	<=	222	;
						10'd168	:	dt	<=	175	;
						10'd169	:	dt	<=	179	;
						10'd170	:	dt	<=	185	;
						10'd171	:	dt	<=	189	;
						10'd172	:	dt	<=	194	;
						10'd173	:	dt	<=	198	;
						10'd174	:	dt	<=	201	;
						10'd175	:	dt	<=	203	;
						10'd176	:	dt	<=	206	;
						10'd177	:	dt	<=	211	;
						10'd178	:	dt	<=	212	;
						10'd179	:	dt	<=	217	;
						10'd180	:	dt	<=	226	;
						10'd181	:	dt	<=	186	;
						10'd182	:	dt	<=	169	;
						10'd183	:	dt	<=	180	;
						10'd184	:	dt	<=	229	;
						10'd185	:	dt	<=	203	;
						10'd186	:	dt	<=	151	;
						10'd187	:	dt	<=	119	;
						10'd188	:	dt	<=	175	;
						10'd189	:	dt	<=	153	;
						10'd190	:	dt	<=	133	;
						10'd191	:	dt	<=	226	;
						10'd192	:	dt	<=	224	;
						10'd193	:	dt	<=	223	;
						10'd194	:	dt	<=	222	;
						10'd195	:	dt	<=	222	;
						10'd196	:	dt	<=	177	;
						10'd197	:	dt	<=	180	;
						10'd198	:	dt	<=	186	;
						10'd199	:	dt	<=	190	;
						10'd200	:	dt	<=	196	;
						10'd201	:	dt	<=	199	;
						10'd202	:	dt	<=	201	;
						10'd203	:	dt	<=	206	;
						10'd204	:	dt	<=	208	;
						10'd205	:	dt	<=	212	;
						10'd206	:	dt	<=	203	;
						10'd207	:	dt	<=	236	;
						10'd208	:	dt	<=	250	;
						10'd209	:	dt	<=	217	;
						10'd210	:	dt	<=	181	;
						10'd211	:	dt	<=	140	;
						10'd212	:	dt	<=	193	;
						10'd213	:	dt	<=	232	;
						10'd214	:	dt	<=	178	;
						10'd215	:	dt	<=	122	;
						10'd216	:	dt	<=	180	;
						10'd217	:	dt	<=	151	;
						10'd218	:	dt	<=	132	;
						10'd219	:	dt	<=	225	;
						10'd220	:	dt	<=	225	;
						10'd221	:	dt	<=	224	;
						10'd222	:	dt	<=	224	;
						10'd223	:	dt	<=	223	;
						10'd224	:	dt	<=	177	;
						10'd225	:	dt	<=	180	;
						10'd226	:	dt	<=	188	;
						10'd227	:	dt	<=	192	;
						10'd228	:	dt	<=	197	;
						10'd229	:	dt	<=	200	;
						10'd230	:	dt	<=	203	;
						10'd231	:	dt	<=	206	;
						10'd232	:	dt	<=	209	;
						10'd233	:	dt	<=	225	;
						10'd234	:	dt	<=	180	;
						10'd235	:	dt	<=	164	;
						10'd236	:	dt	<=	239	;
						10'd237	:	dt	<=	244	;
						10'd238	:	dt	<=	207	;
						10'd239	:	dt	<=	146	;
						10'd240	:	dt	<=	126	;
						10'd241	:	dt	<=	229	;
						10'd242	:	dt	<=	183	;
						10'd243	:	dt	<=	123	;
						10'd244	:	dt	<=	186	;
						10'd245	:	dt	<=	162	;
						10'd246	:	dt	<=	142	;
						10'd247	:	dt	<=	231	;
						10'd248	:	dt	<=	224	;
						10'd249	:	dt	<=	226	;
						10'd250	:	dt	<=	225	;
						10'd251	:	dt	<=	225	;
						10'd252	:	dt	<=	179	;
						10'd253	:	dt	<=	183	;
						10'd254	:	dt	<=	188	;
						10'd255	:	dt	<=	193	;
						10'd256	:	dt	<=	198	;
						10'd257	:	dt	<=	201	;
						10'd258	:	dt	<=	204	;
						10'd259	:	dt	<=	205	;
						10'd260	:	dt	<=	235	;
						10'd261	:	dt	<=	241	;
						10'd262	:	dt	<=	197	;
						10'd263	:	dt	<=	143	;
						10'd264	:	dt	<=	163	;
						10'd265	:	dt	<=	255	;
						10'd266	:	dt	<=	221	;
						10'd267	:	dt	<=	168	;
						10'd268	:	dt	<=	100	;
						10'd269	:	dt	<=	143	;
						10'd270	:	dt	<=	166	;
						10'd271	:	dt	<=	113	;
						10'd272	:	dt	<=	212	;
						10'd273	:	dt	<=	168	;
						10'd274	:	dt	<=	173	;
						10'd275	:	dt	<=	234	;
						10'd276	:	dt	<=	225	;
						10'd277	:	dt	<=	227	;
						10'd278	:	dt	<=	226	;
						10'd279	:	dt	<=	225	;
						10'd280	:	dt	<=	181	;
						10'd281	:	dt	<=	184	;
						10'd282	:	dt	<=	189	;
						10'd283	:	dt	<=	195	;
						10'd284	:	dt	<=	199	;
						10'd285	:	dt	<=	203	;
						10'd286	:	dt	<=	202	;
						10'd287	:	dt	<=	231	;
						10'd288	:	dt	<=	233	;
						10'd289	:	dt	<=	239	;
						10'd290	:	dt	<=	223	;
						10'd291	:	dt	<=	175	;
						10'd292	:	dt	<=	112	;
						10'd293	:	dt	<=	224	;
						10'd294	:	dt	<=	215	;
						10'd295	:	dt	<=	161	;
						10'd296	:	dt	<=	105	;
						10'd297	:	dt	<=	86	;
						10'd298	:	dt	<=	113	;
						10'd299	:	dt	<=	114	;
						10'd300	:	dt	<=	188	;
						10'd301	:	dt	<=	146	;
						10'd302	:	dt	<=	192	;
						10'd303	:	dt	<=	237	;
						10'd304	:	dt	<=	226	;
						10'd305	:	dt	<=	228	;
						10'd306	:	dt	<=	227	;
						10'd307	:	dt	<=	226	;
						10'd308	:	dt	<=	181	;
						10'd309	:	dt	<=	185	;
						10'd310	:	dt	<=	192	;
						10'd311	:	dt	<=	197	;
						10'd312	:	dt	<=	201	;
						10'd313	:	dt	<=	201	;
						10'd314	:	dt	<=	218	;
						10'd315	:	dt	<=	238	;
						10'd316	:	dt	<=	190	;
						10'd317	:	dt	<=	217	;
						10'd318	:	dt	<=	230	;
						10'd319	:	dt	<=	186	;
						10'd320	:	dt	<=	108	;
						10'd321	:	dt	<=	181	;
						10'd322	:	dt	<=	208	;
						10'd323	:	dt	<=	150	;
						10'd324	:	dt	<=	104	;
						10'd325	:	dt	<=	82	;
						10'd326	:	dt	<=	122	;
						10'd327	:	dt	<=	159	;
						10'd328	:	dt	<=	171	;
						10'd329	:	dt	<=	147	;
						10'd330	:	dt	<=	148	;
						10'd331	:	dt	<=	233	;
						10'd332	:	dt	<=	230	;
						10'd333	:	dt	<=	229	;
						10'd334	:	dt	<=	229	;
						10'd335	:	dt	<=	228	;
						10'd336	:	dt	<=	183	;
						10'd337	:	dt	<=	187	;
						10'd338	:	dt	<=	195	;
						10'd339	:	dt	<=	199	;
						10'd340	:	dt	<=	202	;
						10'd341	:	dt	<=	204	;
						10'd342	:	dt	<=	243	;
						10'd343	:	dt	<=	237	;
						10'd344	:	dt	<=	197	;
						10'd345	:	dt	<=	198	;
						10'd346	:	dt	<=	210	;
						10'd347	:	dt	<=	166	;
						10'd348	:	dt	<=	110	;
						10'd349	:	dt	<=	152	;
						10'd350	:	dt	<=	206	;
						10'd351	:	dt	<=	169	;
						10'd352	:	dt	<=	101	;
						10'd353	:	dt	<=	113	;
						10'd354	:	dt	<=	182	;
						10'd355	:	dt	<=	189	;
						10'd356	:	dt	<=	164	;
						10'd357	:	dt	<=	149	;
						10'd358	:	dt	<=	134	;
						10'd359	:	dt	<=	194	;
						10'd360	:	dt	<=	239	;
						10'd361	:	dt	<=	228	;
						10'd362	:	dt	<=	231	;
						10'd363	:	dt	<=	229	;
						10'd364	:	dt	<=	186	;
						10'd365	:	dt	<=	190	;
						10'd366	:	dt	<=	196	;
						10'd367	:	dt	<=	201	;
						10'd368	:	dt	<=	202	;
						10'd369	:	dt	<=	216	;
						10'd370	:	dt	<=	237	;
						10'd371	:	dt	<=	212	;
						10'd372	:	dt	<=	177	;
						10'd373	:	dt	<=	180	;
						10'd374	:	dt	<=	194	;
						10'd375	:	dt	<=	146	;
						10'd376	:	dt	<=	98	;
						10'd377	:	dt	<=	126	;
						10'd378	:	dt	<=	218	;
						10'd379	:	dt	<=	181	;
						10'd380	:	dt	<=	107	;
						10'd381	:	dt	<=	185	;
						10'd382	:	dt	<=	216	;
						10'd383	:	dt	<=	193	;
						10'd384	:	dt	<=	160	;
						10'd385	:	dt	<=	135	;
						10'd386	:	dt	<=	140	;
						10'd387	:	dt	<=	150	;
						10'd388	:	dt	<=	237	;
						10'd389	:	dt	<=	230	;
						10'd390	:	dt	<=	231	;
						10'd391	:	dt	<=	231	;
						10'd392	:	dt	<=	187	;
						10'd393	:	dt	<=	192	;
						10'd394	:	dt	<=	199	;
						10'd395	:	dt	<=	205	;
						10'd396	:	dt	<=	204	;
						10'd397	:	dt	<=	227	;
						10'd398	:	dt	<=	247	;
						10'd399	:	dt	<=	219	;
						10'd400	:	dt	<=	185	;
						10'd401	:	dt	<=	161	;
						10'd402	:	dt	<=	177	;
						10'd403	:	dt	<=	147	;
						10'd404	:	dt	<=	95	;
						10'd405	:	dt	<=	89	;
						10'd406	:	dt	<=	203	;
						10'd407	:	dt	<=	166	;
						10'd408	:	dt	<=	154	;
						10'd409	:	dt	<=	230	;
						10'd410	:	dt	<=	212	;
						10'd411	:	dt	<=	187	;
						10'd412	:	dt	<=	159	;
						10'd413	:	dt	<=	139	;
						10'd414	:	dt	<=	128	;
						10'd415	:	dt	<=	145	;
						10'd416	:	dt	<=	238	;
						10'd417	:	dt	<=	232	;
						10'd418	:	dt	<=	232	;
						10'd419	:	dt	<=	232	;
						10'd420	:	dt	<=	188	;
						10'd421	:	dt	<=	194	;
						10'd422	:	dt	<=	202	;
						10'd423	:	dt	<=	208	;
						10'd424	:	dt	<=	206	;
						10'd425	:	dt	<=	231	;
						10'd426	:	dt	<=	251	;
						10'd427	:	dt	<=	223	;
						10'd428	:	dt	<=	199	;
						10'd429	:	dt	<=	153	;
						10'd430	:	dt	<=	149	;
						10'd431	:	dt	<=	140	;
						10'd432	:	dt	<=	97	;
						10'd433	:	dt	<=	130	;
						10'd434	:	dt	<=	210	;
						10'd435	:	dt	<=	210	;
						10'd436	:	dt	<=	227	;
						10'd437	:	dt	<=	221	;
						10'd438	:	dt	<=	199	;
						10'd439	:	dt	<=	172	;
						10'd440	:	dt	<=	154	;
						10'd441	:	dt	<=	135	;
						10'd442	:	dt	<=	110	;
						10'd443	:	dt	<=	187	;
						10'd444	:	dt	<=	243	;
						10'd445	:	dt	<=	232	;
						10'd446	:	dt	<=	235	;
						10'd447	:	dt	<=	234	;
						10'd448	:	dt	<=	189	;
						10'd449	:	dt	<=	196	;
						10'd450	:	dt	<=	204	;
						10'd451	:	dt	<=	210	;
						10'd452	:	dt	<=	208	;
						10'd453	:	dt	<=	238	;
						10'd454	:	dt	<=	255	;
						10'd455	:	dt	<=	232	;
						10'd456	:	dt	<=	205	;
						10'd457	:	dt	<=	167	;
						10'd458	:	dt	<=	143	;
						10'd459	:	dt	<=	146	;
						10'd460	:	dt	<=	173	;
						10'd461	:	dt	<=	215	;
						10'd462	:	dt	<=	238	;
						10'd463	:	dt	<=	241	;
						10'd464	:	dt	<=	234	;
						10'd465	:	dt	<=	211	;
						10'd466	:	dt	<=	187	;
						10'd467	:	dt	<=	163	;
						10'd468	:	dt	<=	147	;
						10'd469	:	dt	<=	124	;
						10'd470	:	dt	<=	124	;
						10'd471	:	dt	<=	231	;
						10'd472	:	dt	<=	236	;
						10'd473	:	dt	<=	235	;
						10'd474	:	dt	<=	235	;
						10'd475	:	dt	<=	234	;
						10'd476	:	dt	<=	190	;
						10'd477	:	dt	<=	198	;
						10'd478	:	dt	<=	206	;
						10'd479	:	dt	<=	212	;
						10'd480	:	dt	<=	210	;
						10'd481	:	dt	<=	243	;
						10'd482	:	dt	<=	255	;
						10'd483	:	dt	<=	241	;
						10'd484	:	dt	<=	205	;
						10'd485	:	dt	<=	184	;
						10'd486	:	dt	<=	192	;
						10'd487	:	dt	<=	186	;
						10'd488	:	dt	<=	199	;
						10'd489	:	dt	<=	220	;
						10'd490	:	dt	<=	235	;
						10'd491	:	dt	<=	231	;
						10'd492	:	dt	<=	225	;
						10'd493	:	dt	<=	202	;
						10'd494	:	dt	<=	177	;
						10'd495	:	dt	<=	160	;
						10'd496	:	dt	<=	139	;
						10'd497	:	dt	<=	108	;
						10'd498	:	dt	<=	158	;
						10'd499	:	dt	<=	247	;
						10'd500	:	dt	<=	233	;
						10'd501	:	dt	<=	236	;
						10'd502	:	dt	<=	236	;
						10'd503	:	dt	<=	236	;
						10'd504	:	dt	<=	194	;
						10'd505	:	dt	<=	202	;
						10'd506	:	dt	<=	210	;
						10'd507	:	dt	<=	215	;
						10'd508	:	dt	<=	214	;
						10'd509	:	dt	<=	245	;
						10'd510	:	dt	<=	252	;
						10'd511	:	dt	<=	249	;
						10'd512	:	dt	<=	215	;
						10'd513	:	dt	<=	201	;
						10'd514	:	dt	<=	203	;
						10'd515	:	dt	<=	179	;
						10'd516	:	dt	<=	212	;
						10'd517	:	dt	<=	223	;
						10'd518	:	dt	<=	231	;
						10'd519	:	dt	<=	232	;
						10'd520	:	dt	<=	213	;
						10'd521	:	dt	<=	190	;
						10'd522	:	dt	<=	170	;
						10'd523	:	dt	<=	151	;
						10'd524	:	dt	<=	132	;
						10'd525	:	dt	<=	100	;
						10'd526	:	dt	<=	197	;
						10'd527	:	dt	<=	246	;
						10'd528	:	dt	<=	236	;
						10'd529	:	dt	<=	237	;
						10'd530	:	dt	<=	237	;
						10'd531	:	dt	<=	237	;
						10'd532	:	dt	<=	198	;
						10'd533	:	dt	<=	206	;
						10'd534	:	dt	<=	213	;
						10'd535	:	dt	<=	219	;
						10'd536	:	dt	<=	219	;
						10'd537	:	dt	<=	236	;
						10'd538	:	dt	<=	247	;
						10'd539	:	dt	<=	253	;
						10'd540	:	dt	<=	228	;
						10'd541	:	dt	<=	213	;
						10'd542	:	dt	<=	205	;
						10'd543	:	dt	<=	188	;
						10'd544	:	dt	<=	216	;
						10'd545	:	dt	<=	234	;
						10'd546	:	dt	<=	222	;
						10'd547	:	dt	<=	218	;
						10'd548	:	dt	<=	196	;
						10'd549	:	dt	<=	176	;
						10'd550	:	dt	<=	158	;
						10'd551	:	dt	<=	144	;
						10'd552	:	dt	<=	114	;
						10'd553	:	dt	<=	129	;
						10'd554	:	dt	<=	244	;
						10'd555	:	dt	<=	240	;
						10'd556	:	dt	<=	240	;
						10'd557	:	dt	<=	239	;
						10'd558	:	dt	<=	239	;
						10'd559	:	dt	<=	239	;
						10'd560	:	dt	<=	200	;
						10'd561	:	dt	<=	208	;
						10'd562	:	dt	<=	216	;
						10'd563	:	dt	<=	221	;
						10'd564	:	dt	<=	223	;
						10'd565	:	dt	<=	226	;
						10'd566	:	dt	<=	248	;
						10'd567	:	dt	<=	248	;
						10'd568	:	dt	<=	236	;
						10'd569	:	dt	<=	218	;
						10'd570	:	dt	<=	204	;
						10'd571	:	dt	<=	193	;
						10'd572	:	dt	<=	208	;
						10'd573	:	dt	<=	229	;
						10'd574	:	dt	<=	219	;
						10'd575	:	dt	<=	198	;
						10'd576	:	dt	<=	183	;
						10'd577	:	dt	<=	165	;
						10'd578	:	dt	<=	154	;
						10'd579	:	dt	<=	134	;
						10'd580	:	dt	<=	116	;
						10'd581	:	dt	<=	222	;
						10'd582	:	dt	<=	248	;
						10'd583	:	dt	<=	241	;
						10'd584	:	dt	<=	242	;
						10'd585	:	dt	<=	241	;
						10'd586	:	dt	<=	240	;
						10'd587	:	dt	<=	240	;
						10'd588	:	dt	<=	203	;
						10'd589	:	dt	<=	210	;
						10'd590	:	dt	<=	217	;
						10'd591	:	dt	<=	222	;
						10'd592	:	dt	<=	227	;
						10'd593	:	dt	<=	224	;
						10'd594	:	dt	<=	241	;
						10'd595	:	dt	<=	241	;
						10'd596	:	dt	<=	237	;
						10'd597	:	dt	<=	225	;
						10'd598	:	dt	<=	215	;
						10'd599	:	dt	<=	203	;
						10'd600	:	dt	<=	200	;
						10'd601	:	dt	<=	220	;
						10'd602	:	dt	<=	215	;
						10'd603	:	dt	<=	191	;
						10'd604	:	dt	<=	172	;
						10'd605	:	dt	<=	155	;
						10'd606	:	dt	<=	148	;
						10'd607	:	dt	<=	116	;
						10'd608	:	dt	<=	199	;
						10'd609	:	dt	<=	255	;
						10'd610	:	dt	<=	242	;
						10'd611	:	dt	<=	244	;
						10'd612	:	dt	<=	243	;
						10'd613	:	dt	<=	243	;
						10'd614	:	dt	<=	240	;
						10'd615	:	dt	<=	240	;
						10'd616	:	dt	<=	205	;
						10'd617	:	dt	<=	213	;
						10'd618	:	dt	<=	219	;
						10'd619	:	dt	<=	223	;
						10'd620	:	dt	<=	228	;
						10'd621	:	dt	<=	226	;
						10'd622	:	dt	<=	231	;
						10'd623	:	dt	<=	246	;
						10'd624	:	dt	<=	239	;
						10'd625	:	dt	<=	234	;
						10'd626	:	dt	<=	229	;
						10'd627	:	dt	<=	212	;
						10'd628	:	dt	<=	198	;
						10'd629	:	dt	<=	212	;
						10'd630	:	dt	<=	208	;
						10'd631	:	dt	<=	182	;
						10'd632	:	dt	<=	154	;
						10'd633	:	dt	<=	151	;
						10'd634	:	dt	<=	124	;
						10'd635	:	dt	<=	164	;
						10'd636	:	dt	<=	255	;
						10'd637	:	dt	<=	244	;
						10'd638	:	dt	<=	246	;
						10'd639	:	dt	<=	247	;
						10'd640	:	dt	<=	244	;
						10'd641	:	dt	<=	242	;
						10'd642	:	dt	<=	249	;
						10'd643	:	dt	<=	249	;
						10'd644	:	dt	<=	207	;
						10'd645	:	dt	<=	215	;
						10'd646	:	dt	<=	222	;
						10'd647	:	dt	<=	227	;
						10'd648	:	dt	<=	231	;
						10'd649	:	dt	<=	229	;
						10'd650	:	dt	<=	225	;
						10'd651	:	dt	<=	247	;
						10'd652	:	dt	<=	233	;
						10'd653	:	dt	<=	228	;
						10'd654	:	dt	<=	223	;
						10'd655	:	dt	<=	205	;
						10'd656	:	dt	<=	192	;
						10'd657	:	dt	<=	201	;
						10'd658	:	dt	<=	193	;
						10'd659	:	dt	<=	171	;
						10'd660	:	dt	<=	143	;
						10'd661	:	dt	<=	140	;
						10'd662	:	dt	<=	131	;
						10'd663	:	dt	<=	238	;
						10'd664	:	dt	<=	250	;
						10'd665	:	dt	<=	247	;
						10'd666	:	dt	<=	248	;
						10'd667	:	dt	<=	247	;
						10'd668	:	dt	<=	246	;
						10'd669	:	dt	<=	252	;
						10'd670	:	dt	<=	220	;
						10'd671	:	dt	<=	168	;
						10'd672	:	dt	<=	208	;
						10'd673	:	dt	<=	217	;
						10'd674	:	dt	<=	225	;
						10'd675	:	dt	<=	230	;
						10'd676	:	dt	<=	232	;
						10'd677	:	dt	<=	232	;
						10'd678	:	dt	<=	228	;
						10'd679	:	dt	<=	241	;
						10'd680	:	dt	<=	210	;
						10'd681	:	dt	<=	210	;
						10'd682	:	dt	<=	217	;
						10'd683	:	dt	<=	207	;
						10'd684	:	dt	<=	194	;
						10'd685	:	dt	<=	195	;
						10'd686	:	dt	<=	183	;
						10'd687	:	dt	<=	166	;
						10'd688	:	dt	<=	149	;
						10'd689	:	dt	<=	120	;
						10'd690	:	dt	<=	187	;
						10'd691	:	dt	<=	255	;
						10'd692	:	dt	<=	248	;
						10'd693	:	dt	<=	250	;
						10'd694	:	dt	<=	248	;
						10'd695	:	dt	<=	250	;
						10'd696	:	dt	<=	255	;
						10'd697	:	dt	<=	187	;
						10'd698	:	dt	<=	107	;
						10'd699	:	dt	<=	86	;
						10'd700	:	dt	<=	210	;
						10'd701	:	dt	<=	218	;
						10'd702	:	dt	<=	226	;
						10'd703	:	dt	<=	230	;
						10'd704	:	dt	<=	234	;
						10'd705	:	dt	<=	234	;
						10'd706	:	dt	<=	229	;
						10'd707	:	dt	<=	248	;
						10'd708	:	dt	<=	217	;
						10'd709	:	dt	<=	220	;
						10'd710	:	dt	<=	227	;
						10'd711	:	dt	<=	220	;
						10'd712	:	dt	<=	197	;
						10'd713	:	dt	<=	185	;
						10'd714	:	dt	<=	178	;
						10'd715	:	dt	<=	167	;
						10'd716	:	dt	<=	149	;
						10'd717	:	dt	<=	118	;
						10'd718	:	dt	<=	222	;
						10'd719	:	dt	<=	253	;
						10'd720	:	dt	<=	252	;
						10'd721	:	dt	<=	251	;
						10'd722	:	dt	<=	255	;
						10'd723	:	dt	<=	255	;
						10'd724	:	dt	<=	178	;
						10'd725	:	dt	<=	100	;
						10'd726	:	dt	<=	100	;
						10'd727	:	dt	<=	79	;
						10'd728	:	dt	<=	210	;
						10'd729	:	dt	<=	220	;
						10'd730	:	dt	<=	225	;
						10'd731	:	dt	<=	229	;
						10'd732	:	dt	<=	233	;
						10'd733	:	dt	<=	235	;
						10'd734	:	dt	<=	225	;
						10'd735	:	dt	<=	252	;
						10'd736	:	dt	<=	228	;
						10'd737	:	dt	<=	231	;
						10'd738	:	dt	<=	237	;
						10'd739	:	dt	<=	220	;
						10'd740	:	dt	<=	202	;
						10'd741	:	dt	<=	181	;
						10'd742	:	dt	<=	177	;
						10'd743	:	dt	<=	166	;
						10'd744	:	dt	<=	147	;
						10'd745	:	dt	<=	121	;
						10'd746	:	dt	<=	237	;
						10'd747	:	dt	<=	253	;
						10'd748	:	dt	<=	252	;
						10'd749	:	dt	<=	255	;
						10'd750	:	dt	<=	212	;
						10'd751	:	dt	<=	141	;
						10'd752	:	dt	<=	94	;
						10'd753	:	dt	<=	101	;
						10'd754	:	dt	<=	110	;
						10'd755	:	dt	<=	80	;
						10'd756	:	dt	<=	211	;
						10'd757	:	dt	<=	221	;
						10'd758	:	dt	<=	227	;
						10'd759	:	dt	<=	231	;
						10'd760	:	dt	<=	233	;
						10'd761	:	dt	<=	238	;
						10'd762	:	dt	<=	227	;
						10'd763	:	dt	<=	248	;
						10'd764	:	dt	<=	245	;
						10'd765	:	dt	<=	246	;
						10'd766	:	dt	<=	244	;
						10'd767	:	dt	<=	222	;
						10'd768	:	dt	<=	205	;
						10'd769	:	dt	<=	184	;
						10'd770	:	dt	<=	175	;
						10'd771	:	dt	<=	167	;
						10'd772	:	dt	<=	143	;
						10'd773	:	dt	<=	123	;
						10'd774	:	dt	<=	241	;
						10'd775	:	dt	<=	251	;
						10'd776	:	dt	<=	255	;
						10'd777	:	dt	<=	212	;
						10'd778	:	dt	<=	111	;
						10'd779	:	dt	<=	93	;
						10'd780	:	dt	<=	81	;
						10'd781	:	dt	<=	91	;
						10'd782	:	dt	<=	109	;
						10'd783	:	dt	<=	96	;	
					endcase
				end
				5'd14	:	begin
					case (cnt)
						10'd0	:	dt	<=	177	;
						10'd1	:	dt	<=	177	;
						10'd2	:	dt	<=	177	;
						10'd3	:	dt	<=	177	;
						10'd4	:	dt	<=	177	;
						10'd5	:	dt	<=	178	;
						10'd6	:	dt	<=	179	;
						10'd7	:	dt	<=	179	;
						10'd8	:	dt	<=	178	;
						10'd9	:	dt	<=	179	;
						10'd10	:	dt	<=	179	;
						10'd11	:	dt	<=	178	;
						10'd12	:	dt	<=	179	;
						10'd13	:	dt	<=	178	;
						10'd14	:	dt	<=	179	;
						10'd15	:	dt	<=	179	;
						10'd16	:	dt	<=	179	;
						10'd17	:	dt	<=	179	;
						10'd18	:	dt	<=	178	;
						10'd19	:	dt	<=	178	;
						10'd20	:	dt	<=	179	;
						10'd21	:	dt	<=	178	;
						10'd22	:	dt	<=	177	;
						10'd23	:	dt	<=	178	;
						10'd24	:	dt	<=	177	;
						10'd25	:	dt	<=	177	;
						10'd26	:	dt	<=	179	;
						10'd27	:	dt	<=	143	;
						10'd28	:	dt	<=	180	;
						10'd29	:	dt	<=	180	;
						10'd30	:	dt	<=	180	;
						10'd31	:	dt	<=	180	;
						10'd32	:	dt	<=	180	;
						10'd33	:	dt	<=	180	;
						10'd34	:	dt	<=	181	;
						10'd35	:	dt	<=	182	;
						10'd36	:	dt	<=	183	;
						10'd37	:	dt	<=	182	;
						10'd38	:	dt	<=	183	;
						10'd39	:	dt	<=	182	;
						10'd40	:	dt	<=	181	;
						10'd41	:	dt	<=	181	;
						10'd42	:	dt	<=	181	;
						10'd43	:	dt	<=	181	;
						10'd44	:	dt	<=	182	;
						10'd45	:	dt	<=	183	;
						10'd46	:	dt	<=	181	;
						10'd47	:	dt	<=	181	;
						10'd48	:	dt	<=	181	;
						10'd49	:	dt	<=	180	;
						10'd50	:	dt	<=	179	;
						10'd51	:	dt	<=	180	;
						10'd52	:	dt	<=	179	;
						10'd53	:	dt	<=	177	;
						10'd54	:	dt	<=	182	;
						10'd55	:	dt	<=	127	;
						10'd56	:	dt	<=	182	;
						10'd57	:	dt	<=	182	;
						10'd58	:	dt	<=	182	;
						10'd59	:	dt	<=	181	;
						10'd60	:	dt	<=	183	;
						10'd61	:	dt	<=	183	;
						10'd62	:	dt	<=	183	;
						10'd63	:	dt	<=	184	;
						10'd64	:	dt	<=	183	;
						10'd65	:	dt	<=	183	;
						10'd66	:	dt	<=	182	;
						10'd67	:	dt	<=	183	;
						10'd68	:	dt	<=	183	;
						10'd69	:	dt	<=	184	;
						10'd70	:	dt	<=	182	;
						10'd71	:	dt	<=	186	;
						10'd72	:	dt	<=	187	;
						10'd73	:	dt	<=	183	;
						10'd74	:	dt	<=	184	;
						10'd75	:	dt	<=	184	;
						10'd76	:	dt	<=	184	;
						10'd77	:	dt	<=	182	;
						10'd78	:	dt	<=	181	;
						10'd79	:	dt	<=	181	;
						10'd80	:	dt	<=	180	;
						10'd81	:	dt	<=	181	;
						10'd82	:	dt	<=	182	;
						10'd83	:	dt	<=	157	;
						10'd84	:	dt	<=	185	;
						10'd85	:	dt	<=	184	;
						10'd86	:	dt	<=	184	;
						10'd87	:	dt	<=	186	;
						10'd88	:	dt	<=	186	;
						10'd89	:	dt	<=	186	;
						10'd90	:	dt	<=	185	;
						10'd91	:	dt	<=	185	;
						10'd92	:	dt	<=	188	;
						10'd93	:	dt	<=	193	;
						10'd94	:	dt	<=	183	;
						10'd95	:	dt	<=	173	;
						10'd96	:	dt	<=	186	;
						10'd97	:	dt	<=	185	;
						10'd98	:	dt	<=	172	;
						10'd99	:	dt	<=	169	;
						10'd100	:	dt	<=	182	;
						10'd101	:	dt	<=	188	;
						10'd102	:	dt	<=	188	;
						10'd103	:	dt	<=	186	;
						10'd104	:	dt	<=	186	;
						10'd105	:	dt	<=	186	;
						10'd106	:	dt	<=	185	;
						10'd107	:	dt	<=	185	;
						10'd108	:	dt	<=	183	;
						10'd109	:	dt	<=	183	;
						10'd110	:	dt	<=	183	;
						10'd111	:	dt	<=	174	;
						10'd112	:	dt	<=	188	;
						10'd113	:	dt	<=	188	;
						10'd114	:	dt	<=	188	;
						10'd115	:	dt	<=	190	;
						10'd116	:	dt	<=	189	;
						10'd117	:	dt	<=	188	;
						10'd118	:	dt	<=	186	;
						10'd119	:	dt	<=	197	;
						10'd120	:	dt	<=	211	;
						10'd121	:	dt	<=	178	;
						10'd122	:	dt	<=	173	;
						10'd123	:	dt	<=	171	;
						10'd124	:	dt	<=	174	;
						10'd125	:	dt	<=	162	;
						10'd126	:	dt	<=	134	;
						10'd127	:	dt	<=	149	;
						10'd128	:	dt	<=	166	;
						10'd129	:	dt	<=	171	;
						10'd130	:	dt	<=	176	;
						10'd131	:	dt	<=	192	;
						10'd132	:	dt	<=	188	;
						10'd133	:	dt	<=	190	;
						10'd134	:	dt	<=	190	;
						10'd135	:	dt	<=	188	;
						10'd136	:	dt	<=	186	;
						10'd137	:	dt	<=	185	;
						10'd138	:	dt	<=	186	;
						10'd139	:	dt	<=	182	;
						10'd140	:	dt	<=	191	;
						10'd141	:	dt	<=	191	;
						10'd142	:	dt	<=	190	;
						10'd143	:	dt	<=	193	;
						10'd144	:	dt	<=	190	;
						10'd145	:	dt	<=	197	;
						10'd146	:	dt	<=	209	;
						10'd147	:	dt	<=	205	;
						10'd148	:	dt	<=	188	;
						10'd149	:	dt	<=	122	;
						10'd150	:	dt	<=	99	;
						10'd151	:	dt	<=	122	;
						10'd152	:	dt	<=	134	;
						10'd153	:	dt	<=	132	;
						10'd154	:	dt	<=	93	;
						10'd155	:	dt	<=	89	;
						10'd156	:	dt	<=	149	;
						10'd157	:	dt	<=	133	;
						10'd158	:	dt	<=	111	;
						10'd159	:	dt	<=	194	;
						10'd160	:	dt	<=	191	;
						10'd161	:	dt	<=	192	;
						10'd162	:	dt	<=	192	;
						10'd163	:	dt	<=	190	;
						10'd164	:	dt	<=	188	;
						10'd165	:	dt	<=	188	;
						10'd166	:	dt	<=	188	;
						10'd167	:	dt	<=	186	;
						10'd168	:	dt	<=	193	;
						10'd169	:	dt	<=	193	;
						10'd170	:	dt	<=	193	;
						10'd171	:	dt	<=	195	;
						10'd172	:	dt	<=	188	;
						10'd173	:	dt	<=	211	;
						10'd174	:	dt	<=	220	;
						10'd175	:	dt	<=	146	;
						10'd176	:	dt	<=	113	;
						10'd177	:	dt	<=	90	;
						10'd178	:	dt	<=	54	;
						10'd179	:	dt	<=	68	;
						10'd180	:	dt	<=	86	;
						10'd181	:	dt	<=	93	;
						10'd182	:	dt	<=	74	;
						10'd183	:	dt	<=	68	;
						10'd184	:	dt	<=	100	;
						10'd185	:	dt	<=	103	;
						10'd186	:	dt	<=	73	;
						10'd187	:	dt	<=	172	;
						10'd188	:	dt	<=	202	;
						10'd189	:	dt	<=	194	;
						10'd190	:	dt	<=	188	;
						10'd191	:	dt	<=	192	;
						10'd192	:	dt	<=	191	;
						10'd193	:	dt	<=	190	;
						10'd194	:	dt	<=	190	;
						10'd195	:	dt	<=	190	;
						10'd196	:	dt	<=	195	;
						10'd197	:	dt	<=	194	;
						10'd198	:	dt	<=	194	;
						10'd199	:	dt	<=	197	;
						10'd200	:	dt	<=	188	;
						10'd201	:	dt	<=	220	;
						10'd202	:	dt	<=	213	;
						10'd203	:	dt	<=	136	;
						10'd204	:	dt	<=	71	;
						10'd205	:	dt	<=	61	;
						10'd206	:	dt	<=	55	;
						10'd207	:	dt	<=	50	;
						10'd208	:	dt	<=	57	;
						10'd209	:	dt	<=	64	;
						10'd210	:	dt	<=	67	;
						10'd211	:	dt	<=	61	;
						10'd212	:	dt	<=	71	;
						10'd213	:	dt	<=	80	;
						10'd214	:	dt	<=	94	;
						10'd215	:	dt	<=	107	;
						10'd216	:	dt	<=	172	;
						10'd217	:	dt	<=	170	;
						10'd218	:	dt	<=	142	;
						10'd219	:	dt	<=	155	;
						10'd220	:	dt	<=	195	;
						10'd221	:	dt	<=	190	;
						10'd222	:	dt	<=	192	;
						10'd223	:	dt	<=	192	;
						10'd224	:	dt	<=	197	;
						10'd225	:	dt	<=	196	;
						10'd226	:	dt	<=	197	;
						10'd227	:	dt	<=	199	;
						10'd228	:	dt	<=	190	;
						10'd229	:	dt	<=	226	;
						10'd230	:	dt	<=	208	;
						10'd231	:	dt	<=	151	;
						10'd232	:	dt	<=	90	;
						10'd233	:	dt	<=	65	;
						10'd234	:	dt	<=	62	;
						10'd235	:	dt	<=	57	;
						10'd236	:	dt	<=	56	;
						10'd237	:	dt	<=	55	;
						10'd238	:	dt	<=	64	;
						10'd239	:	dt	<=	61	;
						10'd240	:	dt	<=	62	;
						10'd241	:	dt	<=	97	;
						10'd242	:	dt	<=	142	;
						10'd243	:	dt	<=	108	;
						10'd244	:	dt	<=	86	;
						10'd245	:	dt	<=	164	;
						10'd246	:	dt	<=	138	;
						10'd247	:	dt	<=	140	;
						10'd248	:	dt	<=	201	;
						10'd249	:	dt	<=	193	;
						10'd250	:	dt	<=	195	;
						10'd251	:	dt	<=	193	;
						10'd252	:	dt	<=	200	;
						10'd253	:	dt	<=	198	;
						10'd254	:	dt	<=	200	;
						10'd255	:	dt	<=	199	;
						10'd256	:	dt	<=	192	;
						10'd257	:	dt	<=	227	;
						10'd258	:	dt	<=	194	;
						10'd259	:	dt	<=	128	;
						10'd260	:	dt	<=	71	;
						10'd261	:	dt	<=	55	;
						10'd262	:	dt	<=	61	;
						10'd263	:	dt	<=	70	;
						10'd264	:	dt	<=	67	;
						10'd265	:	dt	<=	55	;
						10'd266	:	dt	<=	65	;
						10'd267	:	dt	<=	69	;
						10'd268	:	dt	<=	64	;
						10'd269	:	dt	<=	78	;
						10'd270	:	dt	<=	97	;
						10'd271	:	dt	<=	71	;
						10'd272	:	dt	<=	136	;
						10'd273	:	dt	<=	185	;
						10'd274	:	dt	<=	110	;
						10'd275	:	dt	<=	164	;
						10'd276	:	dt	<=	205	;
						10'd277	:	dt	<=	196	;
						10'd278	:	dt	<=	197	;
						10'd279	:	dt	<=	196	;
						10'd280	:	dt	<=	200	;
						10'd281	:	dt	<=	199	;
						10'd282	:	dt	<=	201	;
						10'd283	:	dt	<=	199	;
						10'd284	:	dt	<=	203	;
						10'd285	:	dt	<=	228	;
						10'd286	:	dt	<=	191	;
						10'd287	:	dt	<=	148	;
						10'd288	:	dt	<=	104	;
						10'd289	:	dt	<=	68	;
						10'd290	:	dt	<=	55	;
						10'd291	:	dt	<=	67	;
						10'd292	:	dt	<=	59	;
						10'd293	:	dt	<=	71	;
						10'd294	:	dt	<=	63	;
						10'd295	:	dt	<=	86	;
						10'd296	:	dt	<=	138	;
						10'd297	:	dt	<=	173	;
						10'd298	:	dt	<=	151	;
						10'd299	:	dt	<=	120	;
						10'd300	:	dt	<=	185	;
						10'd301	:	dt	<=	172	;
						10'd302	:	dt	<=	100	;
						10'd303	:	dt	<=	175	;
						10'd304	:	dt	<=	206	;
						10'd305	:	dt	<=	198	;
						10'd306	:	dt	<=	198	;
						10'd307	:	dt	<=	198	;
						10'd308	:	dt	<=	202	;
						10'd309	:	dt	<=	202	;
						10'd310	:	dt	<=	203	;
						10'd311	:	dt	<=	200	;
						10'd312	:	dt	<=	211	;
						10'd313	:	dt	<=	231	;
						10'd314	:	dt	<=	198	;
						10'd315	:	dt	<=	162	;
						10'd316	:	dt	<=	127	;
						10'd317	:	dt	<=	93	;
						10'd318	:	dt	<=	78	;
						10'd319	:	dt	<=	59	;
						10'd320	:	dt	<=	62	;
						10'd321	:	dt	<=	94	;
						10'd322	:	dt	<=	72	;
						10'd323	:	dt	<=	135	;
						10'd324	:	dt	<=	220	;
						10'd325	:	dt	<=	205	;
						10'd326	:	dt	<=	213	;
						10'd327	:	dt	<=	191	;
						10'd328	:	dt	<=	189	;
						10'd329	:	dt	<=	170	;
						10'd330	:	dt	<=	98	;
						10'd331	:	dt	<=	169	;
						10'd332	:	dt	<=	208	;
						10'd333	:	dt	<=	199	;
						10'd334	:	dt	<=	200	;
						10'd335	:	dt	<=	200	;
						10'd336	:	dt	<=	205	;
						10'd337	:	dt	<=	205	;
						10'd338	:	dt	<=	206	;
						10'd339	:	dt	<=	200	;
						10'd340	:	dt	<=	218	;
						10'd341	:	dt	<=	237	;
						10'd342	:	dt	<=	207	;
						10'd343	:	dt	<=	167	;
						10'd344	:	dt	<=	115	;
						10'd345	:	dt	<=	90	;
						10'd346	:	dt	<=	82	;
						10'd347	:	dt	<=	76	;
						10'd348	:	dt	<=	76	;
						10'd349	:	dt	<=	80	;
						10'd350	:	dt	<=	74	;
						10'd351	:	dt	<=	175	;
						10'd352	:	dt	<=	211	;
						10'd353	:	dt	<=	202	;
						10'd354	:	dt	<=	204	;
						10'd355	:	dt	<=	177	;
						10'd356	:	dt	<=	185	;
						10'd357	:	dt	<=	161	;
						10'd358	:	dt	<=	99	;
						10'd359	:	dt	<=	158	;
						10'd360	:	dt	<=	212	;
						10'd361	:	dt	<=	200	;
						10'd362	:	dt	<=	201	;
						10'd363	:	dt	<=	201	;
						10'd364	:	dt	<=	205	;
						10'd365	:	dt	<=	206	;
						10'd366	:	dt	<=	207	;
						10'd367	:	dt	<=	201	;
						10'd368	:	dt	<=	221	;
						10'd369	:	dt	<=	243	;
						10'd370	:	dt	<=	213	;
						10'd371	:	dt	<=	168	;
						10'd372	:	dt	<=	108	;
						10'd373	:	dt	<=	83	;
						10'd374	:	dt	<=	77	;
						10'd375	:	dt	<=	74	;
						10'd376	:	dt	<=	91	;
						10'd377	:	dt	<=	76	;
						10'd378	:	dt	<=	97	;
						10'd379	:	dt	<=	212	;
						10'd380	:	dt	<=	205	;
						10'd381	:	dt	<=	208	;
						10'd382	:	dt	<=	197	;
						10'd383	:	dt	<=	183	;
						10'd384	:	dt	<=	187	;
						10'd385	:	dt	<=	156	;
						10'd386	:	dt	<=	98	;
						10'd387	:	dt	<=	135	;
						10'd388	:	dt	<=	216	;
						10'd389	:	dt	<=	202	;
						10'd390	:	dt	<=	202	;
						10'd391	:	dt	<=	202	;
						10'd392	:	dt	<=	206	;
						10'd393	:	dt	<=	207	;
						10'd394	:	dt	<=	207	;
						10'd395	:	dt	<=	204	;
						10'd396	:	dt	<=	222	;
						10'd397	:	dt	<=	242	;
						10'd398	:	dt	<=	215	;
						10'd399	:	dt	<=	181	;
						10'd400	:	dt	<=	131	;
						10'd401	:	dt	<=	89	;
						10'd402	:	dt	<=	69	;
						10'd403	:	dt	<=	70	;
						10'd404	:	dt	<=	88	;
						10'd405	:	dt	<=	74	;
						10'd406	:	dt	<=	129	;
						10'd407	:	dt	<=	222	;
						10'd408	:	dt	<=	203	;
						10'd409	:	dt	<=	209	;
						10'd410	:	dt	<=	187	;
						10'd411	:	dt	<=	199	;
						10'd412	:	dt	<=	191	;
						10'd413	:	dt	<=	149	;
						10'd414	:	dt	<=	86	;
						10'd415	:	dt	<=	163	;
						10'd416	:	dt	<=	215	;
						10'd417	:	dt	<=	203	;
						10'd418	:	dt	<=	205	;
						10'd419	:	dt	<=	204	;
						10'd420	:	dt	<=	206	;
						10'd421	:	dt	<=	207	;
						10'd422	:	dt	<=	210	;
						10'd423	:	dt	<=	203	;
						10'd424	:	dt	<=	220	;
						10'd425	:	dt	<=	245	;
						10'd426	:	dt	<=	218	;
						10'd427	:	dt	<=	183	;
						10'd428	:	dt	<=	144	;
						10'd429	:	dt	<=	101	;
						10'd430	:	dt	<=	70	;
						10'd431	:	dt	<=	68	;
						10'd432	:	dt	<=	81	;
						10'd433	:	dt	<=	63	;
						10'd434	:	dt	<=	147	;
						10'd435	:	dt	<=	212	;
						10'd436	:	dt	<=	211	;
						10'd437	:	dt	<=	200	;
						10'd438	:	dt	<=	176	;
						10'd439	:	dt	<=	201	;
						10'd440	:	dt	<=	192	;
						10'd441	:	dt	<=	125	;
						10'd442	:	dt	<=	110	;
						10'd443	:	dt	<=	214	;
						10'd444	:	dt	<=	208	;
						10'd445	:	dt	<=	207	;
						10'd446	:	dt	<=	207	;
						10'd447	:	dt	<=	206	;
						10'd448	:	dt	<=	209	;
						10'd449	:	dt	<=	210	;
						10'd450	:	dt	<=	213	;
						10'd451	:	dt	<=	201	;
						10'd452	:	dt	<=	214	;
						10'd453	:	dt	<=	244	;
						10'd454	:	dt	<=	220	;
						10'd455	:	dt	<=	191	;
						10'd456	:	dt	<=	154	;
						10'd457	:	dt	<=	106	;
						10'd458	:	dt	<=	77	;
						10'd459	:	dt	<=	72	;
						10'd460	:	dt	<=	69	;
						10'd461	:	dt	<=	67	;
						10'd462	:	dt	<=	109	;
						10'd463	:	dt	<=	130	;
						10'd464	:	dt	<=	171	;
						10'd465	:	dt	<=	169	;
						10'd466	:	dt	<=	178	;
						10'd467	:	dt	<=	191	;
						10'd468	:	dt	<=	173	;
						10'd469	:	dt	<=	102	;
						10'd470	:	dt	<=	171	;
						10'd471	:	dt	<=	219	;
						10'd472	:	dt	<=	207	;
						10'd473	:	dt	<=	210	;
						10'd474	:	dt	<=	207	;
						10'd475	:	dt	<=	207	;
						10'd476	:	dt	<=	211	;
						10'd477	:	dt	<=	211	;
						10'd478	:	dt	<=	213	;
						10'd479	:	dt	<=	202	;
						10'd480	:	dt	<=	214	;
						10'd481	:	dt	<=	243	;
						10'd482	:	dt	<=	221	;
						10'd483	:	dt	<=	193	;
						10'd484	:	dt	<=	162	;
						10'd485	:	dt	<=	121	;
						10'd486	:	dt	<=	86	;
						10'd487	:	dt	<=	57	;
						10'd488	:	dt	<=	72	;
						10'd489	:	dt	<=	84	;
						10'd490	:	dt	<=	100	;
						10'd491	:	dt	<=	128	;
						10'd492	:	dt	<=	146	;
						10'd493	:	dt	<=	156	;
						10'd494	:	dt	<=	173	;
						10'd495	:	dt	<=	177	;
						10'd496	:	dt	<=	139	;
						10'd497	:	dt	<=	113	;
						10'd498	:	dt	<=	211	;
						10'd499	:	dt	<=	211	;
						10'd500	:	dt	<=	212	;
						10'd501	:	dt	<=	213	;
						10'd502	:	dt	<=	211	;
						10'd503	:	dt	<=	209	;
						10'd504	:	dt	<=	211	;
						10'd505	:	dt	<=	211	;
						10'd506	:	dt	<=	214	;
						10'd507	:	dt	<=	204	;
						10'd508	:	dt	<=	215	;
						10'd509	:	dt	<=	242	;
						10'd510	:	dt	<=	226	;
						10'd511	:	dt	<=	196	;
						10'd512	:	dt	<=	167	;
						10'd513	:	dt	<=	133	;
						10'd514	:	dt	<=	100	;
						10'd515	:	dt	<=	59	;
						10'd516	:	dt	<=	77	;
						10'd517	:	dt	<=	90	;
						10'd518	:	dt	<=	120	;
						10'd519	:	dt	<=	148	;
						10'd520	:	dt	<=	159	;
						10'd521	:	dt	<=	155	;
						10'd522	:	dt	<=	150	;
						10'd523	:	dt	<=	150	;
						10'd524	:	dt	<=	106	;
						10'd525	:	dt	<=	158	;
						10'd526	:	dt	<=	222	;
						10'd527	:	dt	<=	212	;
						10'd528	:	dt	<=	214	;
						10'd529	:	dt	<=	214	;
						10'd530	:	dt	<=	212	;
						10'd531	:	dt	<=	210	;
						10'd532	:	dt	<=	213	;
						10'd533	:	dt	<=	212	;
						10'd534	:	dt	<=	215	;
						10'd535	:	dt	<=	203	;
						10'd536	:	dt	<=	213	;
						10'd537	:	dt	<=	241	;
						10'd538	:	dt	<=	227	;
						10'd539	:	dt	<=	201	;
						10'd540	:	dt	<=	172	;
						10'd541	:	dt	<=	138	;
						10'd542	:	dt	<=	108	;
						10'd543	:	dt	<=	72	;
						10'd544	:	dt	<=	76	;
						10'd545	:	dt	<=	104	;
						10'd546	:	dt	<=	139	;
						10'd547	:	dt	<=	161	;
						10'd548	:	dt	<=	164	;
						10'd549	:	dt	<=	144	;
						10'd550	:	dt	<=	130	;
						10'd551	:	dt	<=	114	;
						10'd552	:	dt	<=	94	;
						10'd553	:	dt	<=	204	;
						10'd554	:	dt	<=	217	;
						10'd555	:	dt	<=	215	;
						10'd556	:	dt	<=	214	;
						10'd557	:	dt	<=	214	;
						10'd558	:	dt	<=	213	;
						10'd559	:	dt	<=	213	;
						10'd560	:	dt	<=	214	;
						10'd561	:	dt	<=	212	;
						10'd562	:	dt	<=	216	;
						10'd563	:	dt	<=	203	;
						10'd564	:	dt	<=	206	;
						10'd565	:	dt	<=	240	;
						10'd566	:	dt	<=	225	;
						10'd567	:	dt	<=	205	;
						10'd568	:	dt	<=	175	;
						10'd569	:	dt	<=	143	;
						10'd570	:	dt	<=	111	;
						10'd571	:	dt	<=	87	;
						10'd572	:	dt	<=	75	;
						10'd573	:	dt	<=	103	;
						10'd574	:	dt	<=	142	;
						10'd575	:	dt	<=	161	;
						10'd576	:	dt	<=	161	;
						10'd577	:	dt	<=	141	;
						10'd578	:	dt	<=	112	;
						10'd579	:	dt	<=	93	;
						10'd580	:	dt	<=	121	;
						10'd581	:	dt	<=	225	;
						10'd582	:	dt	<=	212	;
						10'd583	:	dt	<=	214	;
						10'd584	:	dt	<=	214	;
						10'd585	:	dt	<=	215	;
						10'd586	:	dt	<=	216	;
						10'd587	:	dt	<=	215	;
						10'd588	:	dt	<=	215	;
						10'd589	:	dt	<=	213	;
						10'd590	:	dt	<=	217	;
						10'd591	:	dt	<=	206	;
						10'd592	:	dt	<=	204	;
						10'd593	:	dt	<=	236	;
						10'd594	:	dt	<=	225	;
						10'd595	:	dt	<=	208	;
						10'd596	:	dt	<=	179	;
						10'd597	:	dt	<=	150	;
						10'd598	:	dt	<=	115	;
						10'd599	:	dt	<=	97	;
						10'd600	:	dt	<=	77	;
						10'd601	:	dt	<=	94	;
						10'd602	:	dt	<=	139	;
						10'd603	:	dt	<=	160	;
						10'd604	:	dt	<=	155	;
						10'd605	:	dt	<=	127	;
						10'd606	:	dt	<=	102	;
						10'd607	:	dt	<=	95	;
						10'd608	:	dt	<=	192	;
						10'd609	:	dt	<=	221	;
						10'd610	:	dt	<=	216	;
						10'd611	:	dt	<=	216	;
						10'd612	:	dt	<=	215	;
						10'd613	:	dt	<=	215	;
						10'd614	:	dt	<=	215	;
						10'd615	:	dt	<=	214	;
						10'd616	:	dt	<=	217	;
						10'd617	:	dt	<=	217	;
						10'd618	:	dt	<=	217	;
						10'd619	:	dt	<=	205	;
						10'd620	:	dt	<=	208	;
						10'd621	:	dt	<=	233	;
						10'd622	:	dt	<=	225	;
						10'd623	:	dt	<=	209	;
						10'd624	:	dt	<=	183	;
						10'd625	:	dt	<=	157	;
						10'd626	:	dt	<=	123	;
						10'd627	:	dt	<=	106	;
						10'd628	:	dt	<=	89	;
						10'd629	:	dt	<=	90	;
						10'd630	:	dt	<=	145	;
						10'd631	:	dt	<=	157	;
						10'd632	:	dt	<=	145	;
						10'd633	:	dt	<=	118	;
						10'd634	:	dt	<=	85	;
						10'd635	:	dt	<=	144	;
						10'd636	:	dt	<=	231	;
						10'd637	:	dt	<=	216	;
						10'd638	:	dt	<=	218	;
						10'd639	:	dt	<=	217	;
						10'd640	:	dt	<=	216	;
						10'd641	:	dt	<=	216	;
						10'd642	:	dt	<=	216	;
						10'd643	:	dt	<=	215	;
						10'd644	:	dt	<=	219	;
						10'd645	:	dt	<=	218	;
						10'd646	:	dt	<=	220	;
						10'd647	:	dt	<=	203	;
						10'd648	:	dt	<=	212	;
						10'd649	:	dt	<=	238	;
						10'd650	:	dt	<=	224	;
						10'd651	:	dt	<=	207	;
						10'd652	:	dt	<=	189	;
						10'd653	:	dt	<=	164	;
						10'd654	:	dt	<=	123	;
						10'd655	:	dt	<=	111	;
						10'd656	:	dt	<=	104	;
						10'd657	:	dt	<=	85	;
						10'd658	:	dt	<=	142	;
						10'd659	:	dt	<=	142	;
						10'd660	:	dt	<=	128	;
						10'd661	:	dt	<=	109	;
						10'd662	:	dt	<=	80	;
						10'd663	:	dt	<=	191	;
						10'd664	:	dt	<=	227	;
						10'd665	:	dt	<=	218	;
						10'd666	:	dt	<=	219	;
						10'd667	:	dt	<=	219	;
						10'd668	:	dt	<=	217	;
						10'd669	:	dt	<=	217	;
						10'd670	:	dt	<=	218	;
						10'd671	:	dt	<=	217	;
						10'd672	:	dt	<=	219	;
						10'd673	:	dt	<=	219	;
						10'd674	:	dt	<=	224	;
						10'd675	:	dt	<=	204	;
						10'd676	:	dt	<=	218	;
						10'd677	:	dt	<=	241	;
						10'd678	:	dt	<=	221	;
						10'd679	:	dt	<=	207	;
						10'd680	:	dt	<=	195	;
						10'd681	:	dt	<=	168	;
						10'd682	:	dt	<=	127	;
						10'd683	:	dt	<=	112	;
						10'd684	:	dt	<=	107	;
						10'd685	:	dt	<=	88	;
						10'd686	:	dt	<=	122	;
						10'd687	:	dt	<=	128	;
						10'd688	:	dt	<=	121	;
						10'd689	:	dt	<=	96	;
						10'd690	:	dt	<=	104	;
						10'd691	:	dt	<=	224	;
						10'd692	:	dt	<=	222	;
						10'd693	:	dt	<=	220	;
						10'd694	:	dt	<=	219	;
						10'd695	:	dt	<=	219	;
						10'd696	:	dt	<=	219	;
						10'd697	:	dt	<=	218	;
						10'd698	:	dt	<=	218	;
						10'd699	:	dt	<=	217	;
						10'd700	:	dt	<=	220	;
						10'd701	:	dt	<=	219	;
						10'd702	:	dt	<=	222	;
						10'd703	:	dt	<=	205	;
						10'd704	:	dt	<=	231	;
						10'd705	:	dt	<=	237	;
						10'd706	:	dt	<=	224	;
						10'd707	:	dt	<=	219	;
						10'd708	:	dt	<=	196	;
						10'd709	:	dt	<=	169	;
						10'd710	:	dt	<=	128	;
						10'd711	:	dt	<=	111	;
						10'd712	:	dt	<=	103	;
						10'd713	:	dt	<=	92	;
						10'd714	:	dt	<=	108	;
						10'd715	:	dt	<=	115	;
						10'd716	:	dt	<=	112	;
						10'd717	:	dt	<=	80	;
						10'd718	:	dt	<=	166	;
						10'd719	:	dt	<=	233	;
						10'd720	:	dt	<=	222	;
						10'd721	:	dt	<=	222	;
						10'd722	:	dt	<=	221	;
						10'd723	:	dt	<=	220	;
						10'd724	:	dt	<=	219	;
						10'd725	:	dt	<=	218	;
						10'd726	:	dt	<=	218	;
						10'd727	:	dt	<=	218	;
						10'd728	:	dt	<=	220	;
						10'd729	:	dt	<=	220	;
						10'd730	:	dt	<=	216	;
						10'd731	:	dt	<=	204	;
						10'd732	:	dt	<=	239	;
						10'd733	:	dt	<=	238	;
						10'd734	:	dt	<=	227	;
						10'd735	:	dt	<=	214	;
						10'd736	:	dt	<=	187	;
						10'd737	:	dt	<=	154	;
						10'd738	:	dt	<=	121	;
						10'd739	:	dt	<=	106	;
						10'd740	:	dt	<=	99	;
						10'd741	:	dt	<=	94	;
						10'd742	:	dt	<=	101	;
						10'd743	:	dt	<=	103	;
						10'd744	:	dt	<=	92	;
						10'd745	:	dt	<=	118	;
						10'd746	:	dt	<=	225	;
						10'd747	:	dt	<=	225	;
						10'd748	:	dt	<=	223	;
						10'd749	:	dt	<=	223	;
						10'd750	:	dt	<=	222	;
						10'd751	:	dt	<=	220	;
						10'd752	:	dt	<=	220	;
						10'd753	:	dt	<=	220	;
						10'd754	:	dt	<=	219	;
						10'd755	:	dt	<=	219	;
						10'd756	:	dt	<=	221	;
						10'd757	:	dt	<=	222	;
						10'd758	:	dt	<=	209	;
						10'd759	:	dt	<=	205	;
						10'd760	:	dt	<=	234	;
						10'd761	:	dt	<=	235	;
						10'd762	:	dt	<=	224	;
						10'd763	:	dt	<=	199	;
						10'd764	:	dt	<=	167	;
						10'd765	:	dt	<=	137	;
						10'd766	:	dt	<=	113	;
						10'd767	:	dt	<=	100	;
						10'd768	:	dt	<=	94	;
						10'd769	:	dt	<=	98	;
						10'd770	:	dt	<=	100	;
						10'd771	:	dt	<=	100	;
						10'd772	:	dt	<=	94	;
						10'd773	:	dt	<=	198	;
						10'd774	:	dt	<=	232	;
						10'd775	:	dt	<=	223	;
						10'd776	:	dt	<=	224	;
						10'd777	:	dt	<=	224	;
						10'd778	:	dt	<=	223	;
						10'd779	:	dt	<=	221	;
						10'd780	:	dt	<=	221	;
						10'd781	:	dt	<=	221	;
						10'd782	:	dt	<=	220	;
						10'd783	:	dt	<=	219	;
					endcase
				end
				5'd15	:	begin
					case (cnt)
						10'd0	:	dt	<=	204	;
						10'd1	:	dt	<=	178	;
						10'd2	:	dt	<=	181	;
						10'd3	:	dt	<=	161	;
						10'd4	:	dt	<=	119	;
						10'd5	:	dt	<=	203	;
						10'd6	:	dt	<=	98	;
						10'd7	:	dt	<=	48	;
						10'd8	:	dt	<=	109	;
						10'd9	:	dt	<=	107	;
						10'd10	:	dt	<=	109	;
						10'd11	:	dt	<=	113	;
						10'd12	:	dt	<=	118	;
						10'd13	:	dt	<=	120	;
						10'd14	:	dt	<=	133	;
						10'd15	:	dt	<=	147	;
						10'd16	:	dt	<=	162	;
						10'd17	:	dt	<=	174	;
						10'd18	:	dt	<=	178	;
						10'd19	:	dt	<=	181	;
						10'd20	:	dt	<=	189	;
						10'd21	:	dt	<=	197	;
						10'd22	:	dt	<=	201	;
						10'd23	:	dt	<=	205	;
						10'd24	:	dt	<=	208	;
						10'd25	:	dt	<=	212	;
						10'd26	:	dt	<=	216	;
						10'd27	:	dt	<=	219	;
						10'd28	:	dt	<=	204	;
						10'd29	:	dt	<=	179	;
						10'd30	:	dt	<=	188	;
						10'd31	:	dt	<=	153	;
						10'd32	:	dt	<=	131	;
						10'd33	:	dt	<=	207	;
						10'd34	:	dt	<=	82	;
						10'd35	:	dt	<=	56	;
						10'd36	:	dt	<=	111	;
						10'd37	:	dt	<=	108	;
						10'd38	:	dt	<=	111	;
						10'd39	:	dt	<=	113	;
						10'd40	:	dt	<=	117	;
						10'd41	:	dt	<=	120	;
						10'd42	:	dt	<=	134	;
						10'd43	:	dt	<=	150	;
						10'd44	:	dt	<=	165	;
						10'd45	:	dt	<=	176	;
						10'd46	:	dt	<=	179	;
						10'd47	:	dt	<=	185	;
						10'd48	:	dt	<=	192	;
						10'd49	:	dt	<=	199	;
						10'd50	:	dt	<=	205	;
						10'd51	:	dt	<=	208	;
						10'd52	:	dt	<=	212	;
						10'd53	:	dt	<=	215	;
						10'd54	:	dt	<=	218	;
						10'd55	:	dt	<=	221	;
						10'd56	:	dt	<=	205	;
						10'd57	:	dt	<=	184	;
						10'd58	:	dt	<=	196	;
						10'd59	:	dt	<=	144	;
						10'd60	:	dt	<=	147	;
						10'd61	:	dt	<=	207	;
						10'd62	:	dt	<=	68	;
						10'd63	:	dt	<=	68	;
						10'd64	:	dt	<=	113	;
						10'd65	:	dt	<=	108	;
						10'd66	:	dt	<=	112	;
						10'd67	:	dt	<=	116	;
						10'd68	:	dt	<=	119	;
						10'd69	:	dt	<=	120	;
						10'd70	:	dt	<=	136	;
						10'd71	:	dt	<=	153	;
						10'd72	:	dt	<=	167	;
						10'd73	:	dt	<=	178	;
						10'd74	:	dt	<=	183	;
						10'd75	:	dt	<=	187	;
						10'd76	:	dt	<=	194	;
						10'd77	:	dt	<=	202	;
						10'd78	:	dt	<=	207	;
						10'd79	:	dt	<=	210	;
						10'd80	:	dt	<=	215	;
						10'd81	:	dt	<=	218	;
						10'd82	:	dt	<=	221	;
						10'd83	:	dt	<=	225	;
						10'd84	:	dt	<=	202	;
						10'd85	:	dt	<=	187	;
						10'd86	:	dt	<=	200	;
						10'd87	:	dt	<=	137	;
						10'd88	:	dt	<=	163	;
						10'd89	:	dt	<=	200	;
						10'd90	:	dt	<=	57	;
						10'd91	:	dt	<=	80	;
						10'd92	:	dt	<=	114	;
						10'd93	:	dt	<=	109	;
						10'd94	:	dt	<=	113	;
						10'd95	:	dt	<=	116	;
						10'd96	:	dt	<=	118	;
						10'd97	:	dt	<=	123	;
						10'd98	:	dt	<=	139	;
						10'd99	:	dt	<=	155	;
						10'd100	:	dt	<=	170	;
						10'd101	:	dt	<=	181	;
						10'd102	:	dt	<=	184	;
						10'd103	:	dt	<=	189	;
						10'd104	:	dt	<=	197	;
						10'd105	:	dt	<=	205	;
						10'd106	:	dt	<=	211	;
						10'd107	:	dt	<=	215	;
						10'd108	:	dt	<=	218	;
						10'd109	:	dt	<=	222	;
						10'd110	:	dt	<=	225	;
						10'd111	:	dt	<=	227	;
						10'd112	:	dt	<=	202	;
						10'd113	:	dt	<=	188	;
						10'd114	:	dt	<=	201	;
						10'd115	:	dt	<=	126	;
						10'd116	:	dt	<=	182	;
						10'd117	:	dt	<=	189	;
						10'd118	:	dt	<=	39	;
						10'd119	:	dt	<=	86	;
						10'd120	:	dt	<=	111	;
						10'd121	:	dt	<=	107	;
						10'd122	:	dt	<=	112	;
						10'd123	:	dt	<=	118	;
						10'd124	:	dt	<=	124	;
						10'd125	:	dt	<=	125	;
						10'd126	:	dt	<=	143	;
						10'd127	:	dt	<=	162	;
						10'd128	:	dt	<=	175	;
						10'd129	:	dt	<=	185	;
						10'd130	:	dt	<=	187	;
						10'd131	:	dt	<=	191	;
						10'd132	:	dt	<=	201	;
						10'd133	:	dt	<=	209	;
						10'd134	:	dt	<=	213	;
						10'd135	:	dt	<=	218	;
						10'd136	:	dt	<=	222	;
						10'd137	:	dt	<=	226	;
						10'd138	:	dt	<=	229	;
						10'd139	:	dt	<=	231	;
						10'd140	:	dt	<=	198	;
						10'd141	:	dt	<=	200	;
						10'd142	:	dt	<=	196	;
						10'd143	:	dt	<=	144	;
						10'd144	:	dt	<=	180	;
						10'd145	:	dt	<=	174	;
						10'd146	:	dt	<=	115	;
						10'd147	:	dt	<=	136	;
						10'd148	:	dt	<=	137	;
						10'd149	:	dt	<=	144	;
						10'd150	:	dt	<=	154	;
						10'd151	:	dt	<=	156	;
						10'd152	:	dt	<=	153	;
						10'd153	:	dt	<=	131	;
						10'd154	:	dt	<=	132	;
						10'd155	:	dt	<=	147	;
						10'd156	:	dt	<=	163	;
						10'd157	:	dt	<=	181	;
						10'd158	:	dt	<=	190	;
						10'd159	:	dt	<=	196	;
						10'd160	:	dt	<=	204	;
						10'd161	:	dt	<=	212	;
						10'd162	:	dt	<=	224	;
						10'd163	:	dt	<=	227	;
						10'd164	:	dt	<=	224	;
						10'd165	:	dt	<=	229	;
						10'd166	:	dt	<=	232	;
						10'd167	:	dt	<=	236	;
						10'd168	:	dt	<=	194	;
						10'd169	:	dt	<=	214	;
						10'd170	:	dt	<=	181	;
						10'd171	:	dt	<=	158	;
						10'd172	:	dt	<=	159	;
						10'd173	:	dt	<=	157	;
						10'd174	:	dt	<=	159	;
						10'd175	:	dt	<=	145	;
						10'd176	:	dt	<=	137	;
						10'd177	:	dt	<=	145	;
						10'd178	:	dt	<=	141	;
						10'd179	:	dt	<=	136	;
						10'd180	:	dt	<=	128	;
						10'd181	:	dt	<=	137	;
						10'd182	:	dt	<=	136	;
						10'd183	:	dt	<=	133	;
						10'd184	:	dt	<=	137	;
						10'd185	:	dt	<=	143	;
						10'd186	:	dt	<=	154	;
						10'd187	:	dt	<=	165	;
						10'd188	:	dt	<=	165	;
						10'd189	:	dt	<=	159	;
						10'd190	:	dt	<=	173	;
						10'd191	:	dt	<=	207	;
						10'd192	:	dt	<=	238	;
						10'd193	:	dt	<=	237	;
						10'd194	:	dt	<=	235	;
						10'd195	:	dt	<=	240	;
						10'd196	:	dt	<=	199	;
						10'd197	:	dt	<=	193	;
						10'd198	:	dt	<=	153	;
						10'd199	:	dt	<=	148	;
						10'd200	:	dt	<=	148	;
						10'd201	:	dt	<=	144	;
						10'd202	:	dt	<=	136	;
						10'd203	:	dt	<=	130	;
						10'd204	:	dt	<=	131	;
						10'd205	:	dt	<=	133	;
						10'd206	:	dt	<=	132	;
						10'd207	:	dt	<=	130	;
						10'd208	:	dt	<=	131	;
						10'd209	:	dt	<=	146	;
						10'd210	:	dt	<=	149	;
						10'd211	:	dt	<=	146	;
						10'd212	:	dt	<=	143	;
						10'd213	:	dt	<=	140	;
						10'd214	:	dt	<=	139	;
						10'd215	:	dt	<=	153	;
						10'd216	:	dt	<=	161	;
						10'd217	:	dt	<=	147	;
						10'd218	:	dt	<=	133	;
						10'd219	:	dt	<=	119	;
						10'd220	:	dt	<=	161	;
						10'd221	:	dt	<=	228	;
						10'd222	:	dt	<=	250	;
						10'd223	:	dt	<=	243	;
						10'd224	:	dt	<=	203	;
						10'd225	:	dt	<=	201	;
						10'd226	:	dt	<=	168	;
						10'd227	:	dt	<=	133	;
						10'd228	:	dt	<=	140	;
						10'd229	:	dt	<=	127	;
						10'd230	:	dt	<=	130	;
						10'd231	:	dt	<=	125	;
						10'd232	:	dt	<=	131	;
						10'd233	:	dt	<=	136	;
						10'd234	:	dt	<=	136	;
						10'd235	:	dt	<=	134	;
						10'd236	:	dt	<=	140	;
						10'd237	:	dt	<=	152	;
						10'd238	:	dt	<=	152	;
						10'd239	:	dt	<=	149	;
						10'd240	:	dt	<=	142	;
						10'd241	:	dt	<=	136	;
						10'd242	:	dt	<=	142	;
						10'd243	:	dt	<=	156	;
						10'd244	:	dt	<=	156	;
						10'd245	:	dt	<=	153	;
						10'd246	:	dt	<=	146	;
						10'd247	:	dt	<=	129	;
						10'd248	:	dt	<=	110	;
						10'd249	:	dt	<=	120	;
						10'd250	:	dt	<=	193	;
						10'd251	:	dt	<=	251	;
						10'd252	:	dt	<=	203	;
						10'd253	:	dt	<=	211	;
						10'd254	:	dt	<=	175	;
						10'd255	:	dt	<=	137	;
						10'd256	:	dt	<=	220	;
						10'd257	:	dt	<=	106	;
						10'd258	:	dt	<=	73	;
						10'd259	:	dt	<=	119	;
						10'd260	:	dt	<=	117	;
						10'd261	:	dt	<=	121	;
						10'd262	:	dt	<=	124	;
						10'd263	:	dt	<=	128	;
						10'd264	:	dt	<=	139	;
						10'd265	:	dt	<=	150	;
						10'd266	:	dt	<=	153	;
						10'd267	:	dt	<=	147	;
						10'd268	:	dt	<=	137	;
						10'd269	:	dt	<=	139	;
						10'd270	:	dt	<=	152	;
						10'd271	:	dt	<=	155	;
						10'd272	:	dt	<=	147	;
						10'd273	:	dt	<=	151	;
						10'd274	:	dt	<=	145	;
						10'd275	:	dt	<=	136	;
						10'd276	:	dt	<=	131	;
						10'd277	:	dt	<=	118	;
						10'd278	:	dt	<=	105	;
						10'd279	:	dt	<=	143	;
						10'd280	:	dt	<=	207	;
						10'd281	:	dt	<=	216	;
						10'd282	:	dt	<=	160	;
						10'd283	:	dt	<=	153	;
						10'd284	:	dt	<=	234	;
						10'd285	:	dt	<=	83	;
						10'd286	:	dt	<=	56	;
						10'd287	:	dt	<=	119	;
						10'd288	:	dt	<=	110	;
						10'd289	:	dt	<=	112	;
						10'd290	:	dt	<=	114	;
						10'd291	:	dt	<=	118	;
						10'd292	:	dt	<=	119	;
						10'd293	:	dt	<=	137	;
						10'd294	:	dt	<=	156	;
						10'd295	:	dt	<=	185	;
						10'd296	:	dt	<=	165	;
						10'd297	:	dt	<=	151	;
						10'd298	:	dt	<=	151	;
						10'd299	:	dt	<=	152	;
						10'd300	:	dt	<=	153	;
						10'd301	:	dt	<=	151	;
						10'd302	:	dt	<=	146	;
						10'd303	:	dt	<=	140	;
						10'd304	:	dt	<=	139	;
						10'd305	:	dt	<=	142	;
						10'd306	:	dt	<=	126	;
						10'd307	:	dt	<=	105	;
						10'd308	:	dt	<=	211	;
						10'd309	:	dt	<=	222	;
						10'd310	:	dt	<=	150	;
						10'd311	:	dt	<=	170	;
						10'd312	:	dt	<=	226	;
						10'd313	:	dt	<=	69	;
						10'd314	:	dt	<=	72	;
						10'd315	:	dt	<=	120	;
						10'd316	:	dt	<=	111	;
						10'd317	:	dt	<=	113	;
						10'd318	:	dt	<=	115	;
						10'd319	:	dt	<=	119	;
						10'd320	:	dt	<=	121	;
						10'd321	:	dt	<=	134	;
						10'd322	:	dt	<=	168	;
						10'd323	:	dt	<=	220	;
						10'd324	:	dt	<=	199	;
						10'd325	:	dt	<=	169	;
						10'd326	:	dt	<=	157	;
						10'd327	:	dt	<=	150	;
						10'd328	:	dt	<=	141	;
						10'd329	:	dt	<=	146	;
						10'd330	:	dt	<=	141	;
						10'd331	:	dt	<=	143	;
						10'd332	:	dt	<=	142	;
						10'd333	:	dt	<=	157	;
						10'd334	:	dt	<=	138	;
						10'd335	:	dt	<=	120	;
						10'd336	:	dt	<=	213	;
						10'd337	:	dt	<=	224	;
						10'd338	:	dt	<=	141	;
						10'd339	:	dt	<=	185	;
						10'd340	:	dt	<=	218	;
						10'd341	:	dt	<=	56	;
						10'd342	:	dt	<=	81	;
						10'd343	:	dt	<=	121	;
						10'd344	:	dt	<=	112	;
						10'd345	:	dt	<=	113	;
						10'd346	:	dt	<=	116	;
						10'd347	:	dt	<=	118	;
						10'd348	:	dt	<=	122	;
						10'd349	:	dt	<=	134	;
						10'd350	:	dt	<=	209	;
						10'd351	:	dt	<=	201	;
						10'd352	:	dt	<=	176	;
						10'd353	:	dt	<=	133	;
						10'd354	:	dt	<=	128	;
						10'd355	:	dt	<=	139	;
						10'd356	:	dt	<=	116	;
						10'd357	:	dt	<=	119	;
						10'd358	:	dt	<=	141	;
						10'd359	:	dt	<=	145	;
						10'd360	:	dt	<=	153	;
						10'd361	:	dt	<=	168	;
						10'd362	:	dt	<=	146	;
						10'd363	:	dt	<=	132	;
						10'd364	:	dt	<=	213	;
						10'd365	:	dt	<=	222	;
						10'd366	:	dt	<=	137	;
						10'd367	:	dt	<=	201	;
						10'd368	:	dt	<=	205	;
						10'd369	:	dt	<=	47	;
						10'd370	:	dt	<=	90	;
						10'd371	:	dt	<=	119	;
						10'd372	:	dt	<=	111	;
						10'd373	:	dt	<=	113	;
						10'd374	:	dt	<=	116	;
						10'd375	:	dt	<=	121	;
						10'd376	:	dt	<=	114	;
						10'd377	:	dt	<=	170	;
						10'd378	:	dt	<=	219	;
						10'd379	:	dt	<=	174	;
						10'd380	:	dt	<=	160	;
						10'd381	:	dt	<=	123	;
						10'd382	:	dt	<=	82	;
						10'd383	:	dt	<=	95	;
						10'd384	:	dt	<=	77	;
						10'd385	:	dt	<=	84	;
						10'd386	:	dt	<=	176	;
						10'd387	:	dt	<=	165	;
						10'd388	:	dt	<=	170	;
						10'd389	:	dt	<=	162	;
						10'd390	:	dt	<=	142	;
						10'd391	:	dt	<=	140	;
						10'd392	:	dt	<=	215	;
						10'd393	:	dt	<=	219	;
						10'd394	:	dt	<=	131	;
						10'd395	:	dt	<=	214	;
						10'd396	:	dt	<=	190	;
						10'd397	:	dt	<=	41	;
						10'd398	:	dt	<=	99	;
						10'd399	:	dt	<=	119	;
						10'd400	:	dt	<=	111	;
						10'd401	:	dt	<=	113	;
						10'd402	:	dt	<=	117	;
						10'd403	:	dt	<=	116	;
						10'd404	:	dt	<=	132	;
						10'd405	:	dt	<=	227	;
						10'd406	:	dt	<=	195	;
						10'd407	:	dt	<=	158	;
						10'd408	:	dt	<=	139	;
						10'd409	:	dt	<=	116	;
						10'd410	:	dt	<=	75	;
						10'd411	:	dt	<=	68	;
						10'd412	:	dt	<=	53	;
						10'd413	:	dt	<=	90	;
						10'd414	:	dt	<=	200	;
						10'd415	:	dt	<=	188	;
						10'd416	:	dt	<=	180	;
						10'd417	:	dt	<=	149	;
						10'd418	:	dt	<=	134	;
						10'd419	:	dt	<=	141	;
						10'd420	:	dt	<=	217	;
						10'd421	:	dt	<=	213	;
						10'd422	:	dt	<=	131	;
						10'd423	:	dt	<=	228	;
						10'd424	:	dt	<=	176	;
						10'd425	:	dt	<=	37	;
						10'd426	:	dt	<=	107	;
						10'd427	:	dt	<=	119	;
						10'd428	:	dt	<=	113	;
						10'd429	:	dt	<=	113	;
						10'd430	:	dt	<=	117	;
						10'd431	:	dt	<=	108	;
						10'd432	:	dt	<=	172	;
						10'd433	:	dt	<=	243	;
						10'd434	:	dt	<=	195	;
						10'd435	:	dt	<=	151	;
						10'd436	:	dt	<=	130	;
						10'd437	:	dt	<=	88	;
						10'd438	:	dt	<=	65	;
						10'd439	:	dt	<=	69	;
						10'd440	:	dt	<=	49	;
						10'd441	:	dt	<=	119	;
						10'd442	:	dt	<=	203	;
						10'd443	:	dt	<=	203	;
						10'd444	:	dt	<=	192	;
						10'd445	:	dt	<=	153	;
						10'd446	:	dt	<=	128	;
						10'd447	:	dt	<=	134	;
						10'd448	:	dt	<=	223	;
						10'd449	:	dt	<=	208	;
						10'd450	:	dt	<=	133	;
						10'd451	:	dt	<=	237	;
						10'd452	:	dt	<=	157	;
						10'd453	:	dt	<=	37	;
						10'd454	:	dt	<=	114	;
						10'd455	:	dt	<=	118	;
						10'd456	:	dt	<=	112	;
						10'd457	:	dt	<=	114	;
						10'd458	:	dt	<=	118	;
						10'd459	:	dt	<=	110	;
						10'd460	:	dt	<=	148	;
						10'd461	:	dt	<=	230	;
						10'd462	:	dt	<=	213	;
						10'd463	:	dt	<=	169	;
						10'd464	:	dt	<=	135	;
						10'd465	:	dt	<=	79	;
						10'd466	:	dt	<=	58	;
						10'd467	:	dt	<=	67	;
						10'd468	:	dt	<=	71	;
						10'd469	:	dt	<=	129	;
						10'd470	:	dt	<=	195	;
						10'd471	:	dt	<=	215	;
						10'd472	:	dt	<=	199	;
						10'd473	:	dt	<=	158	;
						10'd474	:	dt	<=	129	;
						10'd475	:	dt	<=	125	;
						10'd476	:	dt	<=	231	;
						10'd477	:	dt	<=	201	;
						10'd478	:	dt	<=	139	;
						10'd479	:	dt	<=	248	;
						10'd480	:	dt	<=	141	;
						10'd481	:	dt	<=	40	;
						10'd482	:	dt	<=	119	;
						10'd483	:	dt	<=	116	;
						10'd484	:	dt	<=	112	;
						10'd485	:	dt	<=	113	;
						10'd486	:	dt	<=	116	;
						10'd487	:	dt	<=	119	;
						10'd488	:	dt	<=	117	;
						10'd489	:	dt	<=	209	;
						10'd490	:	dt	<=	235	;
						10'd491	:	dt	<=	200	;
						10'd492	:	dt	<=	148	;
						10'd493	:	dt	<=	95	;
						10'd494	:	dt	<=	52	;
						10'd495	:	dt	<=	99	;
						10'd496	:	dt	<=	113	;
						10'd497	:	dt	<=	115	;
						10'd498	:	dt	<=	187	;
						10'd499	:	dt	<=	207	;
						10'd500	:	dt	<=	181	;
						10'd501	:	dt	<=	152	;
						10'd502	:	dt	<=	129	;
						10'd503	:	dt	<=	111	;
						10'd504	:	dt	<=	237	;
						10'd505	:	dt	<=	194	;
						10'd506	:	dt	<=	148	;
						10'd507	:	dt	<=	255	;
						10'd508	:	dt	<=	126	;
						10'd509	:	dt	<=	45	;
						10'd510	:	dt	<=	122	;
						10'd511	:	dt	<=	115	;
						10'd512	:	dt	<=	112	;
						10'd513	:	dt	<=	112	;
						10'd514	:	dt	<=	115	;
						10'd515	:	dt	<=	119	;
						10'd516	:	dt	<=	119	;
						10'd517	:	dt	<=	170	;
						10'd518	:	dt	<=	252	;
						10'd519	:	dt	<=	221	;
						10'd520	:	dt	<=	164	;
						10'd521	:	dt	<=	106	;
						10'd522	:	dt	<=	68	;
						10'd523	:	dt	<=	75	;
						10'd524	:	dt	<=	136	;
						10'd525	:	dt	<=	178	;
						10'd526	:	dt	<=	192	;
						10'd527	:	dt	<=	175	;
						10'd528	:	dt	<=	147	;
						10'd529	:	dt	<=	141	;
						10'd530	:	dt	<=	124	;
						10'd531	:	dt	<=	102	;
						10'd532	:	dt	<=	243	;
						10'd533	:	dt	<=	182	;
						10'd534	:	dt	<=	160	;
						10'd535	:	dt	<=	255	;
						10'd536	:	dt	<=	109	;
						10'd537	:	dt	<=	51	;
						10'd538	:	dt	<=	125	;
						10'd539	:	dt	<=	114	;
						10'd540	:	dt	<=	110	;
						10'd541	:	dt	<=	110	;
						10'd542	:	dt	<=	113	;
						10'd543	:	dt	<=	115	;
						10'd544	:	dt	<=	124	;
						10'd545	:	dt	<=	145	;
						10'd546	:	dt	<=	238	;
						10'd547	:	dt	<=	235	;
						10'd548	:	dt	<=	205	;
						10'd549	:	dt	<=	187	;
						10'd550	:	dt	<=	179	;
						10'd551	:	dt	<=	179	;
						10'd552	:	dt	<=	196	;
						10'd553	:	dt	<=	176	;
						10'd554	:	dt	<=	155	;
						10'd555	:	dt	<=	134	;
						10'd556	:	dt	<=	122	;
						10'd557	:	dt	<=	125	;
						10'd558	:	dt	<=	120	;
						10'd559	:	dt	<=	106	;
						10'd560	:	dt	<=	246	;
						10'd561	:	dt	<=	172	;
						10'd562	:	dt	<=	176	;
						10'd563	:	dt	<=	255	;
						10'd564	:	dt	<=	91	;
						10'd565	:	dt	<=	58	;
						10'd566	:	dt	<=	124	;
						10'd567	:	dt	<=	111	;
						10'd568	:	dt	<=	109	;
						10'd569	:	dt	<=	109	;
						10'd570	:	dt	<=	112	;
						10'd571	:	dt	<=	112	;
						10'd572	:	dt	<=	125	;
						10'd573	:	dt	<=	142	;
						10'd574	:	dt	<=	203	;
						10'd575	:	dt	<=	245	;
						10'd576	:	dt	<=	209	;
						10'd577	:	dt	<=	192	;
						10'd578	:	dt	<=	188	;
						10'd579	:	dt	<=	197	;
						10'd580	:	dt	<=	192	;
						10'd581	:	dt	<=	145	;
						10'd582	:	dt	<=	117	;
						10'd583	:	dt	<=	119	;
						10'd584	:	dt	<=	114	;
						10'd585	:	dt	<=	115	;
						10'd586	:	dt	<=	122	;
						10'd587	:	dt	<=	126	;
						10'd588	:	dt	<=	248	;
						10'd589	:	dt	<=	160	;
						10'd590	:	dt	<=	191	;
						10'd591	:	dt	<=	252	;
						10'd592	:	dt	<=	76	;
						10'd593	:	dt	<=	67	;
						10'd594	:	dt	<=	123	;
						10'd595	:	dt	<=	109	;
						10'd596	:	dt	<=	108	;
						10'd597	:	dt	<=	108	;
						10'd598	:	dt	<=	111	;
						10'd599	:	dt	<=	113	;
						10'd600	:	dt	<=	123	;
						10'd601	:	dt	<=	152	;
						10'd602	:	dt	<=	227	;
						10'd603	:	dt	<=	196	;
						10'd604	:	dt	<=	165	;
						10'd605	:	dt	<=	162	;
						10'd606	:	dt	<=	171	;
						10'd607	:	dt	<=	198	;
						10'd608	:	dt	<=	191	;
						10'd609	:	dt	<=	131	;
						10'd610	:	dt	<=	108	;
						10'd611	:	dt	<=	110	;
						10'd612	:	dt	<=	104	;
						10'd613	:	dt	<=	118	;
						10'd614	:	dt	<=	122	;
						10'd615	:	dt	<=	115	;
						10'd616	:	dt	<=	246	;
						10'd617	:	dt	<=	153	;
						10'd618	:	dt	<=	209	;
						10'd619	:	dt	<=	241	;
						10'd620	:	dt	<=	65	;
						10'd621	:	dt	<=	78	;
						10'd622	:	dt	<=	123	;
						10'd623	:	dt	<=	109	;
						10'd624	:	dt	<=	107	;
						10'd625	:	dt	<=	107	;
						10'd626	:	dt	<=	111	;
						10'd627	:	dt	<=	115	;
						10'd628	:	dt	<=	116	;
						10'd629	:	dt	<=	185	;
						10'd630	:	dt	<=	231	;
						10'd631	:	dt	<=	171	;
						10'd632	:	dt	<=	163	;
						10'd633	:	dt	<=	166	;
						10'd634	:	dt	<=	163	;
						10'd635	:	dt	<=	186	;
						10'd636	:	dt	<=	185	;
						10'd637	:	dt	<=	139	;
						10'd638	:	dt	<=	108	;
						10'd639	:	dt	<=	121	;
						10'd640	:	dt	<=	214	;
						10'd641	:	dt	<=	149	;
						10'd642	:	dt	<=	89	;
						10'd643	:	dt	<=	84	;
						10'd644	:	dt	<=	241	;
						10'd645	:	dt	<=	147	;
						10'd646	:	dt	<=	225	;
						10'd647	:	dt	<=	229	;
						10'd648	:	dt	<=	42	;
						10'd649	:	dt	<=	76	;
						10'd650	:	dt	<=	114	;
						10'd651	:	dt	<=	99	;
						10'd652	:	dt	<=	98	;
						10'd653	:	dt	<=	99	;
						10'd654	:	dt	<=	103	;
						10'd655	:	dt	<=	108	;
						10'd656	:	dt	<=	112	;
						10'd657	:	dt	<=	184	;
						10'd658	:	dt	<=	212	;
						10'd659	:	dt	<=	165	;
						10'd660	:	dt	<=	150	;
						10'd661	:	dt	<=	149	;
						10'd662	:	dt	<=	145	;
						10'd663	:	dt	<=	169	;
						10'd664	:	dt	<=	169	;
						10'd665	:	dt	<=	142	;
						10'd666	:	dt	<=	98	;
						10'd667	:	dt	<=	214	;
						10'd668	:	dt	<=	255	;
						10'd669	:	dt	<=	159	;
						10'd670	:	dt	<=	90	;
						10'd671	:	dt	<=	89	;
						10'd672	:	dt	<=	236	;
						10'd673	:	dt	<=	144	;
						10'd674	:	dt	<=	235	;
						10'd675	:	dt	<=	216	;
						10'd676	:	dt	<=	113	;
						10'd677	:	dt	<=	134	;
						10'd678	:	dt	<=	148	;
						10'd679	:	dt	<=	134	;
						10'd680	:	dt	<=	128	;
						10'd681	:	dt	<=	124	;
						10'd682	:	dt	<=	121	;
						10'd683	:	dt	<=	122	;
						10'd684	:	dt	<=	132	;
						10'd685	:	dt	<=	162	;
						10'd686	:	dt	<=	186	;
						10'd687	:	dt	<=	177	;
						10'd688	:	dt	<=	191	;
						10'd689	:	dt	<=	188	;
						10'd690	:	dt	<=	138	;
						10'd691	:	dt	<=	117	;
						10'd692	:	dt	<=	163	;
						10'd693	:	dt	<=	136	;
						10'd694	:	dt	<=	113	;
						10'd695	:	dt	<=	205	;
						10'd696	:	dt	<=	255	;
						10'd697	:	dt	<=	166	;
						10'd698	:	dt	<=	97	;
						10'd699	:	dt	<=	92	;
						10'd700	:	dt	<=	229	;
						10'd701	:	dt	<=	148	;
						10'd702	:	dt	<=	239	;
						10'd703	:	dt	<=	220	;
						10'd704	:	dt	<=	185	;
						10'd705	:	dt	<=	149	;
						10'd706	:	dt	<=	162	;
						10'd707	:	dt	<=	162	;
						10'd708	:	dt	<=	160	;
						10'd709	:	dt	<=	157	;
						10'd710	:	dt	<=	158	;
						10'd711	:	dt	<=	162	;
						10'd712	:	dt	<=	159	;
						10'd713	:	dt	<=	157	;
						10'd714	:	dt	<=	159	;
						10'd715	:	dt	<=	169	;
						10'd716	:	dt	<=	177	;
						10'd717	:	dt	<=	226	;
						10'd718	:	dt	<=	192	;
						10'd719	:	dt	<=	115	;
						10'd720	:	dt	<=	170	;
						10'd721	:	dt	<=	169	;
						10'd722	:	dt	<=	145	;
						10'd723	:	dt	<=	192	;
						10'd724	:	dt	<=	227	;
						10'd725	:	dt	<=	153	;
						10'd726	:	dt	<=	106	;
						10'd727	:	dt	<=	95	;
						10'd728	:	dt	<=	222	;
						10'd729	:	dt	<=	151	;
						10'd730	:	dt	<=	245	;
						10'd731	:	dt	<=	219	;
						10'd732	:	dt	<=	168	;
						10'd733	:	dt	<=	132	;
						10'd734	:	dt	<=	150	;
						10'd735	:	dt	<=	147	;
						10'd736	:	dt	<=	148	;
						10'd737	:	dt	<=	149	;
						10'd738	:	dt	<=	152	;
						10'd739	:	dt	<=	151	;
						10'd740	:	dt	<=	153	;
						10'd741	:	dt	<=	152	;
						10'd742	:	dt	<=	150	;
						10'd743	:	dt	<=	154	;
						10'd744	:	dt	<=	147	;
						10'd745	:	dt	<=	179	;
						10'd746	:	dt	<=	226	;
						10'd747	:	dt	<=	155	;
						10'd748	:	dt	<=	142	;
						10'd749	:	dt	<=	159	;
						10'd750	:	dt	<=	158	;
						10'd751	:	dt	<=	154	;
						10'd752	:	dt	<=	158	;
						10'd753	:	dt	<=	134	;
						10'd754	:	dt	<=	103	;
						10'd755	:	dt	<=	102	;
						10'd756	:	dt	<=	214	;
						10'd757	:	dt	<=	157	;
						10'd758	:	dt	<=	249	;
						10'd759	:	dt	<=	214	;
						10'd760	:	dt	<=	168	;
						10'd761	:	dt	<=	142	;
						10'd762	:	dt	<=	153	;
						10'd763	:	dt	<=	154	;
						10'd764	:	dt	<=	155	;
						10'd765	:	dt	<=	155	;
						10'd766	:	dt	<=	155	;
						10'd767	:	dt	<=	156	;
						10'd768	:	dt	<=	158	;
						10'd769	:	dt	<=	159	;
						10'd770	:	dt	<=	161	;
						10'd771	:	dt	<=	163	;
						10'd772	:	dt	<=	161	;
						10'd773	:	dt	<=	158	;
						10'd774	:	dt	<=	181	;
						10'd775	:	dt	<=	172	;
						10'd776	:	dt	<=	161	;
						10'd777	:	dt	<=	165	;
						10'd778	:	dt	<=	165	;
						10'd779	:	dt	<=	166	;
						10'd780	:	dt	<=	171	;
						10'd781	:	dt	<=	138	;
						10'd782	:	dt	<=	88	;
						10'd783	:	dt	<=	69	;
					endcase
				end
				5'd16	:	begin
					case (cnt)
						10'd0	:	dt	<=	107	;
						10'd1	:	dt	<=	109	;
						10'd2	:	dt	<=	114	;
						10'd3	:	dt	<=	120	;
						10'd4	:	dt	<=	133	;
						10'd5	:	dt	<=	145	;
						10'd6	:	dt	<=	153	;
						10'd7	:	dt	<=	161	;
						10'd8	:	dt	<=	168	;
						10'd9	:	dt	<=	171	;
						10'd10	:	dt	<=	172	;
						10'd11	:	dt	<=	175	;
						10'd12	:	dt	<=	181	;
						10'd13	:	dt	<=	187	;
						10'd14	:	dt	<=	191	;
						10'd15	:	dt	<=	197	;
						10'd16	:	dt	<=	199	;
						10'd17	:	dt	<=	201	;
						10'd18	:	dt	<=	203	;
						10'd19	:	dt	<=	206	;
						10'd20	:	dt	<=	209	;
						10'd21	:	dt	<=	210	;
						10'd22	:	dt	<=	212	;
						10'd23	:	dt	<=	214	;
						10'd24	:	dt	<=	215	;
						10'd25	:	dt	<=	215	;
						10'd26	:	dt	<=	218	;
						10'd27	:	dt	<=	220	;
						10'd28	:	dt	<=	107	;
						10'd29	:	dt	<=	110	;
						10'd30	:	dt	<=	115	;
						10'd31	:	dt	<=	122	;
						10'd32	:	dt	<=	134	;
						10'd33	:	dt	<=	146	;
						10'd34	:	dt	<=	156	;
						10'd35	:	dt	<=	163	;
						10'd36	:	dt	<=	169	;
						10'd37	:	dt	<=	172	;
						10'd38	:	dt	<=	173	;
						10'd39	:	dt	<=	176	;
						10'd40	:	dt	<=	183	;
						10'd41	:	dt	<=	189	;
						10'd42	:	dt	<=	191	;
						10'd43	:	dt	<=	195	;
						10'd44	:	dt	<=	199	;
						10'd45	:	dt	<=	203	;
						10'd46	:	dt	<=	205	;
						10'd47	:	dt	<=	207	;
						10'd48	:	dt	<=	209	;
						10'd49	:	dt	<=	211	;
						10'd50	:	dt	<=	213	;
						10'd51	:	dt	<=	215	;
						10'd52	:	dt	<=	217	;
						10'd53	:	dt	<=	217	;
						10'd54	:	dt	<=	217	;
						10'd55	:	dt	<=	220	;
						10'd56	:	dt	<=	108	;
						10'd57	:	dt	<=	111	;
						10'd58	:	dt	<=	117	;
						10'd59	:	dt	<=	122	;
						10'd60	:	dt	<=	135	;
						10'd61	:	dt	<=	147	;
						10'd62	:	dt	<=	157	;
						10'd63	:	dt	<=	165	;
						10'd64	:	dt	<=	170	;
						10'd65	:	dt	<=	172	;
						10'd66	:	dt	<=	174	;
						10'd67	:	dt	<=	179	;
						10'd68	:	dt	<=	184	;
						10'd69	:	dt	<=	189	;
						10'd70	:	dt	<=	192	;
						10'd71	:	dt	<=	197	;
						10'd72	:	dt	<=	200	;
						10'd73	:	dt	<=	204	;
						10'd74	:	dt	<=	206	;
						10'd75	:	dt	<=	209	;
						10'd76	:	dt	<=	209	;
						10'd77	:	dt	<=	212	;
						10'd78	:	dt	<=	214	;
						10'd79	:	dt	<=	217	;
						10'd80	:	dt	<=	218	;
						10'd81	:	dt	<=	218	;
						10'd82	:	dt	<=	220	;
						10'd83	:	dt	<=	221	;
						10'd84	:	dt	<=	108	;
						10'd85	:	dt	<=	113	;
						10'd86	:	dt	<=	116	;
						10'd87	:	dt	<=	122	;
						10'd88	:	dt	<=	137	;
						10'd89	:	dt	<=	148	;
						10'd90	:	dt	<=	157	;
						10'd91	:	dt	<=	164	;
						10'd92	:	dt	<=	171	;
						10'd93	:	dt	<=	174	;
						10'd94	:	dt	<=	177	;
						10'd95	:	dt	<=	181	;
						10'd96	:	dt	<=	185	;
						10'd97	:	dt	<=	189	;
						10'd98	:	dt	<=	195	;
						10'd99	:	dt	<=	198	;
						10'd100	:	dt	<=	201	;
						10'd101	:	dt	<=	204	;
						10'd102	:	dt	<=	205	;
						10'd103	:	dt	<=	208	;
						10'd104	:	dt	<=	211	;
						10'd105	:	dt	<=	214	;
						10'd106	:	dt	<=	216	;
						10'd107	:	dt	<=	218	;
						10'd108	:	dt	<=	218	;
						10'd109	:	dt	<=	219	;
						10'd110	:	dt	<=	220	;
						10'd111	:	dt	<=	221	;
						10'd112	:	dt	<=	108	;
						10'd113	:	dt	<=	113	;
						10'd114	:	dt	<=	116	;
						10'd115	:	dt	<=	123	;
						10'd116	:	dt	<=	139	;
						10'd117	:	dt	<=	152	;
						10'd118	:	dt	<=	161	;
						10'd119	:	dt	<=	167	;
						10'd120	:	dt	<=	173	;
						10'd121	:	dt	<=	176	;
						10'd122	:	dt	<=	179	;
						10'd123	:	dt	<=	182	;
						10'd124	:	dt	<=	190	;
						10'd125	:	dt	<=	196	;
						10'd126	:	dt	<=	196	;
						10'd127	:	dt	<=	202	;
						10'd128	:	dt	<=	208	;
						10'd129	:	dt	<=	207	;
						10'd130	:	dt	<=	208	;
						10'd131	:	dt	<=	211	;
						10'd132	:	dt	<=	214	;
						10'd133	:	dt	<=	216	;
						10'd134	:	dt	<=	219	;
						10'd135	:	dt	<=	219	;
						10'd136	:	dt	<=	219	;
						10'd137	:	dt	<=	221	;
						10'd138	:	dt	<=	221	;
						10'd139	:	dt	<=	221	;
						10'd140	:	dt	<=	109	;
						10'd141	:	dt	<=	114	;
						10'd142	:	dt	<=	117	;
						10'd143	:	dt	<=	126	;
						10'd144	:	dt	<=	141	;
						10'd145	:	dt	<=	154	;
						10'd146	:	dt	<=	165	;
						10'd147	:	dt	<=	167	;
						10'd148	:	dt	<=	172	;
						10'd149	:	dt	<=	177	;
						10'd150	:	dt	<=	178	;
						10'd151	:	dt	<=	176	;
						10'd152	:	dt	<=	178	;
						10'd153	:	dt	<=	171	;
						10'd154	:	dt	<=	157	;
						10'd155	:	dt	<=	148	;
						10'd156	:	dt	<=	163	;
						10'd157	:	dt	<=	209	;
						10'd158	:	dt	<=	211	;
						10'd159	:	dt	<=	211	;
						10'd160	:	dt	<=	217	;
						10'd161	:	dt	<=	219	;
						10'd162	:	dt	<=	220	;
						10'd163	:	dt	<=	220	;
						10'd164	:	dt	<=	222	;
						10'd165	:	dt	<=	224	;
						10'd166	:	dt	<=	224	;
						10'd167	:	dt	<=	224	;
						10'd168	:	dt	<=	111	;
						10'd169	:	dt	<=	115	;
						10'd170	:	dt	<=	119	;
						10'd171	:	dt	<=	129	;
						10'd172	:	dt	<=	143	;
						10'd173	:	dt	<=	154	;
						10'd174	:	dt	<=	158	;
						10'd175	:	dt	<=	169	;
						10'd176	:	dt	<=	182	;
						10'd177	:	dt	<=	175	;
						10'd178	:	dt	<=	159	;
						10'd179	:	dt	<=	143	;
						10'd180	:	dt	<=	130	;
						10'd181	:	dt	<=	114	;
						10'd182	:	dt	<=	105	;
						10'd183	:	dt	<=	108	;
						10'd184	:	dt	<=	99	;
						10'd185	:	dt	<=	124	;
						10'd186	:	dt	<=	207	;
						10'd187	:	dt	<=	220	;
						10'd188	:	dt	<=	217	;
						10'd189	:	dt	<=	220	;
						10'd190	:	dt	<=	223	;
						10'd191	:	dt	<=	224	;
						10'd192	:	dt	<=	225	;
						10'd193	:	dt	<=	225	;
						10'd194	:	dt	<=	226	;
						10'd195	:	dt	<=	227	;
						10'd196	:	dt	<=	112	;
						10'd197	:	dt	<=	116	;
						10'd198	:	dt	<=	118	;
						10'd199	:	dt	<=	131	;
						10'd200	:	dt	<=	142	;
						10'd201	:	dt	<=	152	;
						10'd202	:	dt	<=	175	;
						10'd203	:	dt	<=	196	;
						10'd204	:	dt	<=	186	;
						10'd205	:	dt	<=	157	;
						10'd206	:	dt	<=	121	;
						10'd207	:	dt	<=	116	;
						10'd208	:	dt	<=	114	;
						10'd209	:	dt	<=	100	;
						10'd210	:	dt	<=	91	;
						10'd211	:	dt	<=	102	;
						10'd212	:	dt	<=	114	;
						10'd213	:	dt	<=	88	;
						10'd214	:	dt	<=	111	;
						10'd215	:	dt	<=	212	;
						10'd216	:	dt	<=	224	;
						10'd217	:	dt	<=	220	;
						10'd218	:	dt	<=	226	;
						10'd219	:	dt	<=	228	;
						10'd220	:	dt	<=	228	;
						10'd221	:	dt	<=	228	;
						10'd222	:	dt	<=	229	;
						10'd223	:	dt	<=	229	;
						10'd224	:	dt	<=	112	;
						10'd225	:	dt	<=	117	;
						10'd226	:	dt	<=	122	;
						10'd227	:	dt	<=	126	;
						10'd228	:	dt	<=	142	;
						10'd229	:	dt	<=	186	;
						10'd230	:	dt	<=	205	;
						10'd231	:	dt	<=	171	;
						10'd232	:	dt	<=	139	;
						10'd233	:	dt	<=	113	;
						10'd234	:	dt	<=	91	;
						10'd235	:	dt	<=	107	;
						10'd236	:	dt	<=	109	;
						10'd237	:	dt	<=	95	;
						10'd238	:	dt	<=	89	;
						10'd239	:	dt	<=	101	;
						10'd240	:	dt	<=	107	;
						10'd241	:	dt	<=	95	;
						10'd242	:	dt	<=	95	;
						10'd243	:	dt	<=	115	;
						10'd244	:	dt	<=	228	;
						10'd245	:	dt	<=	223	;
						10'd246	:	dt	<=	227	;
						10'd247	:	dt	<=	229	;
						10'd248	:	dt	<=	228	;
						10'd249	:	dt	<=	229	;
						10'd250	:	dt	<=	231	;
						10'd251	:	dt	<=	230	;
						10'd252	:	dt	<=	114	;
						10'd253	:	dt	<=	119	;
						10'd254	:	dt	<=	109	;
						10'd255	:	dt	<=	150	;
						10'd256	:	dt	<=	189	;
						10'd257	:	dt	<=	180	;
						10'd258	:	dt	<=	134	;
						10'd259	:	dt	<=	117	;
						10'd260	:	dt	<=	110	;
						10'd261	:	dt	<=	95	;
						10'd262	:	dt	<=	90	;
						10'd263	:	dt	<=	111	;
						10'd264	:	dt	<=	109	;
						10'd265	:	dt	<=	92	;
						10'd266	:	dt	<=	95	;
						10'd267	:	dt	<=	105	;
						10'd268	:	dt	<=	104	;
						10'd269	:	dt	<=	95	;
						10'd270	:	dt	<=	118	;
						10'd271	:	dt	<=	77	;
						10'd272	:	dt	<=	153	;
						10'd273	:	dt	<=	240	;
						10'd274	:	dt	<=	225	;
						10'd275	:	dt	<=	230	;
						10'd276	:	dt	<=	230	;
						10'd277	:	dt	<=	232	;
						10'd278	:	dt	<=	233	;
						10'd279	:	dt	<=	232	;
						10'd280	:	dt	<=	112	;
						10'd281	:	dt	<=	111	;
						10'd282	:	dt	<=	162	;
						10'd283	:	dt	<=	204	;
						10'd284	:	dt	<=	156	;
						10'd285	:	dt	<=	117	;
						10'd286	:	dt	<=	94	;
						10'd287	:	dt	<=	99	;
						10'd288	:	dt	<=	98	;
						10'd289	:	dt	<=	78	;
						10'd290	:	dt	<=	103	;
						10'd291	:	dt	<=	119	;
						10'd292	:	dt	<=	105	;
						10'd293	:	dt	<=	94	;
						10'd294	:	dt	<=	106	;
						10'd295	:	dt	<=	107	;
						10'd296	:	dt	<=	94	;
						10'd297	:	dt	<=	106	;
						10'd298	:	dt	<=	115	;
						10'd299	:	dt	<=	99	;
						10'd300	:	dt	<=	84	;
						10'd301	:	dt	<=	220	;
						10'd302	:	dt	<=	230	;
						10'd303	:	dt	<=	229	;
						10'd304	:	dt	<=	233	;
						10'd305	:	dt	<=	236	;
						10'd306	:	dt	<=	236	;
						10'd307	:	dt	<=	236	;
						10'd308	:	dt	<=	105	;
						10'd309	:	dt	<=	213	;
						10'd310	:	dt	<=	230	;
						10'd311	:	dt	<=	150	;
						10'd312	:	dt	<=	110	;
						10'd313	:	dt	<=	95	;
						10'd314	:	dt	<=	82	;
						10'd315	:	dt	<=	81	;
						10'd316	:	dt	<=	116	;
						10'd317	:	dt	<=	153	;
						10'd318	:	dt	<=	113	;
						10'd319	:	dt	<=	94	;
						10'd320	:	dt	<=	66	;
						10'd321	:	dt	<=	96	;
						10'd322	:	dt	<=	116	;
						10'd323	:	dt	<=	102	;
						10'd324	:	dt	<=	72	;
						10'd325	:	dt	<=	112	;
						10'd326	:	dt	<=	112	;
						10'd327	:	dt	<=	98	;
						10'd328	:	dt	<=	72	;
						10'd329	:	dt	<=	142	;
						10'd330	:	dt	<=	248	;
						10'd331	:	dt	<=	231	;
						10'd332	:	dt	<=	236	;
						10'd333	:	dt	<=	236	;
						10'd334	:	dt	<=	236	;
						10'd335	:	dt	<=	237	;
						10'd336	:	dt	<=	140	;
						10'd337	:	dt	<=	255	;
						10'd338	:	dt	<=	174	;
						10'd339	:	dt	<=	129	;
						10'd340	:	dt	<=	97	;
						10'd341	:	dt	<=	76	;
						10'd342	:	dt	<=	103	;
						10'd343	:	dt	<=	152	;
						10'd344	:	dt	<=	236	;
						10'd345	:	dt	<=	235	;
						10'd346	:	dt	<=	133	;
						10'd347	:	dt	<=	66	;
						10'd348	:	dt	<=	70	;
						10'd349	:	dt	<=	73	;
						10'd350	:	dt	<=	105	;
						10'd351	:	dt	<=	83	;
						10'd352	:	dt	<=	60	;
						10'd353	:	dt	<=	125	;
						10'd354	:	dt	<=	108	;
						10'd355	:	dt	<=	92	;
						10'd356	:	dt	<=	88	;
						10'd357	:	dt	<=	68	;
						10'd358	:	dt	<=	187	;
						10'd359	:	dt	<=	245	;
						10'd360	:	dt	<=	234	;
						10'd361	:	dt	<=	236	;
						10'd362	:	dt	<=	238	;
						10'd363	:	dt	<=	238	;
						10'd364	:	dt	<=	118	;
						10'd365	:	dt	<=	195	;
						10'd366	:	dt	<=	142	;
						10'd367	:	dt	<=	104	;
						10'd368	:	dt	<=	101	;
						10'd369	:	dt	<=	167	;
						10'd370	:	dt	<=	249	;
						10'd371	:	dt	<=	243	;
						10'd372	:	dt	<=	251	;
						10'd373	:	dt	<=	220	;
						10'd374	:	dt	<=	156	;
						10'd375	:	dt	<=	87	;
						10'd376	:	dt	<=	78	;
						10'd377	:	dt	<=	73	;
						10'd378	:	dt	<=	61	;
						10'd379	:	dt	<=	36	;
						10'd380	:	dt	<=	74	;
						10'd381	:	dt	<=	134	;
						10'd382	:	dt	<=	102	;
						10'd383	:	dt	<=	107	;
						10'd384	:	dt	<=	107	;
						10'd385	:	dt	<=	96	;
						10'd386	:	dt	<=	89	;
						10'd387	:	dt	<=	200	;
						10'd388	:	dt	<=	245	;
						10'd389	:	dt	<=	236	;
						10'd390	:	dt	<=	239	;
						10'd391	:	dt	<=	241	;
						10'd392	:	dt	<=	111	;
						10'd393	:	dt	<=	122	;
						10'd394	:	dt	<=	126	;
						10'd395	:	dt	<=	113	;
						10'd396	:	dt	<=	225	;
						10'd397	:	dt	<=	251	;
						10'd398	:	dt	<=	247	;
						10'd399	:	dt	<=	233	;
						10'd400	:	dt	<=	249	;
						10'd401	:	dt	<=	211	;
						10'd402	:	dt	<=	159	;
						10'd403	:	dt	<=	108	;
						10'd404	:	dt	<=	86	;
						10'd405	:	dt	<=	77	;
						10'd406	:	dt	<=	25	;
						10'd407	:	dt	<=	6	;
						10'd408	:	dt	<=	84	;
						10'd409	:	dt	<=	132	;
						10'd410	:	dt	<=	101	;
						10'd411	:	dt	<=	117	;
						10'd412	:	dt	<=	121	;
						10'd413	:	dt	<=	120	;
						10'd414	:	dt	<=	100	;
						10'd415	:	dt	<=	106	;
						10'd416	:	dt	<=	243	;
						10'd417	:	dt	<=	241	;
						10'd418	:	dt	<=	242	;
						10'd419	:	dt	<=	242	;
						10'd420	:	dt	<=	118	;
						10'd421	:	dt	<=	119	;
						10'd422	:	dt	<=	121	;
						10'd423	:	dt	<=	150	;
						10'd424	:	dt	<=	255	;
						10'd425	:	dt	<=	225	;
						10'd426	:	dt	<=	248	;
						10'd427	:	dt	<=	240	;
						10'd428	:	dt	<=	244	;
						10'd429	:	dt	<=	193	;
						10'd430	:	dt	<=	141	;
						10'd431	:	dt	<=	111	;
						10'd432	:	dt	<=	104	;
						10'd433	:	dt	<=	92	;
						10'd434	:	dt	<=	81	;
						10'd435	:	dt	<=	17	;
						10'd436	:	dt	<=	62	;
						10'd437	:	dt	<=	122	;
						10'd438	:	dt	<=	100	;
						10'd439	:	dt	<=	114	;
						10'd440	:	dt	<=	127	;
						10'd441	:	dt	<=	111	;
						10'd442	:	dt	<=	100	;
						10'd443	:	dt	<=	73	;
						10'd444	:	dt	<=	197	;
						10'd445	:	dt	<=	253	;
						10'd446	:	dt	<=	241	;
						10'd447	:	dt	<=	243	;
						10'd448	:	dt	<=	117	;
						10'd449	:	dt	<=	123	;
						10'd450	:	dt	<=	114	;
						10'd451	:	dt	<=	175	;
						10'd452	:	dt	<=	255	;
						10'd453	:	dt	<=	228	;
						10'd454	:	dt	<=	255	;
						10'd455	:	dt	<=	242	;
						10'd456	:	dt	<=	221	;
						10'd457	:	dt	<=	160	;
						10'd458	:	dt	<=	105	;
						10'd459	:	dt	<=	110	;
						10'd460	:	dt	<=	116	;
						10'd461	:	dt	<=	105	;
						10'd462	:	dt	<=	98	;
						10'd463	:	dt	<=	69	;
						10'd464	:	dt	<=	36	;
						10'd465	:	dt	<=	98	;
						10'd466	:	dt	<=	110	;
						10'd467	:	dt	<=	166	;
						10'd468	:	dt	<=	147	;
						10'd469	:	dt	<=	101	;
						10'd470	:	dt	<=	87	;
						10'd471	:	dt	<=	65	;
						10'd472	:	dt	<=	142	;
						10'd473	:	dt	<=	255	;
						10'd474	:	dt	<=	241	;
						10'd475	:	dt	<=	245	;
						10'd476	:	dt	<=	118	;
						10'd477	:	dt	<=	122	;
						10'd478	:	dt	<=	112	;
						10'd479	:	dt	<=	212	;
						10'd480	:	dt	<=	255	;
						10'd481	:	dt	<=	224	;
						10'd482	:	dt	<=	255	;
						10'd483	:	dt	<=	238	;
						10'd484	:	dt	<=	193	;
						10'd485	:	dt	<=	132	;
						10'd486	:	dt	<=	116	;
						10'd487	:	dt	<=	123	;
						10'd488	:	dt	<=	126	;
						10'd489	:	dt	<=	120	;
						10'd490	:	dt	<=	100	;
						10'd491	:	dt	<=	87	;
						10'd492	:	dt	<=	41	;
						10'd493	:	dt	<=	56	;
						10'd494	:	dt	<=	174	;
						10'd495	:	dt	<=	216	;
						10'd496	:	dt	<=	211	;
						10'd497	:	dt	<=	185	;
						10'd498	:	dt	<=	141	;
						10'd499	:	dt	<=	62	;
						10'd500	:	dt	<=	143	;
						10'd501	:	dt	<=	255	;
						10'd502	:	dt	<=	242	;
						10'd503	:	dt	<=	246	;
						10'd504	:	dt	<=	120	;
						10'd505	:	dt	<=	124	;
						10'd506	:	dt	<=	113	;
						10'd507	:	dt	<=	223	;
						10'd508	:	dt	<=	255	;
						10'd509	:	dt	<=	219	;
						10'd510	:	dt	<=	223	;
						10'd511	:	dt	<=	210	;
						10'd512	:	dt	<=	137	;
						10'd513	:	dt	<=	101	;
						10'd514	:	dt	<=	105	;
						10'd515	:	dt	<=	132	;
						10'd516	:	dt	<=	126	;
						10'd517	:	dt	<=	109	;
						10'd518	:	dt	<=	102	;
						10'd519	:	dt	<=	91	;
						10'd520	:	dt	<=	79	;
						10'd521	:	dt	<=	60	;
						10'd522	:	dt	<=	205	;
						10'd523	:	dt	<=	238	;
						10'd524	:	dt	<=	239	;
						10'd525	:	dt	<=	239	;
						10'd526	:	dt	<=	234	;
						10'd527	:	dt	<=	173	;
						10'd528	:	dt	<=	184	;
						10'd529	:	dt	<=	255	;
						10'd530	:	dt	<=	246	;
						10'd531	:	dt	<=	249	;
						10'd532	:	dt	<=	118	;
						10'd533	:	dt	<=	122	;
						10'd534	:	dt	<=	116	;
						10'd535	:	dt	<=	191	;
						10'd536	:	dt	<=	255	;
						10'd537	:	dt	<=	218	;
						10'd538	:	dt	<=	152	;
						10'd539	:	dt	<=	139	;
						10'd540	:	dt	<=	91	;
						10'd541	:	dt	<=	88	;
						10'd542	:	dt	<=	99	;
						10'd543	:	dt	<=	106	;
						10'd544	:	dt	<=	101	;
						10'd545	:	dt	<=	91	;
						10'd546	:	dt	<=	86	;
						10'd547	:	dt	<=	82	;
						10'd548	:	dt	<=	103	;
						10'd549	:	dt	<=	79	;
						10'd550	:	dt	<=	196	;
						10'd551	:	dt	<=	248	;
						10'd552	:	dt	<=	241	;
						10'd553	:	dt	<=	245	;
						10'd554	:	dt	<=	249	;
						10'd555	:	dt	<=	232	;
						10'd556	:	dt	<=	167	;
						10'd557	:	dt	<=	194	;
						10'd558	:	dt	<=	255	;
						10'd559	:	dt	<=	248	;
						10'd560	:	dt	<=	118	;
						10'd561	:	dt	<=	120	;
						10'd562	:	dt	<=	125	;
						10'd563	:	dt	<=	152	;
						10'd564	:	dt	<=	233	;
						10'd565	:	dt	<=	150	;
						10'd566	:	dt	<=	106	;
						10'd567	:	dt	<=	97	;
						10'd568	:	dt	<=	97	;
						10'd569	:	dt	<=	109	;
						10'd570	:	dt	<=	116	;
						10'd571	:	dt	<=	104	;
						10'd572	:	dt	<=	82	;
						10'd573	:	dt	<=	78	;
						10'd574	:	dt	<=	84	;
						10'd575	:	dt	<=	75	;
						10'd576	:	dt	<=	82	;
						10'd577	:	dt	<=	66	;
						10'd578	:	dt	<=	157	;
						10'd579	:	dt	<=	255	;
						10'd580	:	dt	<=	233	;
						10'd581	:	dt	<=	241	;
						10'd582	:	dt	<=	241	;
						10'd583	:	dt	<=	210	;
						10'd584	:	dt	<=	155	;
						10'd585	:	dt	<=	128	;
						10'd586	:	dt	<=	255	;
						10'd587	:	dt	<=	249	;
						10'd588	:	dt	<=	119	;
						10'd589	:	dt	<=	119	;
						10'd590	:	dt	<=	129	;
						10'd591	:	dt	<=	143	;
						10'd592	:	dt	<=	171	;
						10'd593	:	dt	<=	116	;
						10'd594	:	dt	<=	95	;
						10'd595	:	dt	<=	117	;
						10'd596	:	dt	<=	110	;
						10'd597	:	dt	<=	93	;
						10'd598	:	dt	<=	84	;
						10'd599	:	dt	<=	79	;
						10'd600	:	dt	<=	69	;
						10'd601	:	dt	<=	65	;
						10'd602	:	dt	<=	69	;
						10'd603	:	dt	<=	65	;
						10'd604	:	dt	<=	83	;
						10'd605	:	dt	<=	107	;
						10'd606	:	dt	<=	115	;
						10'd607	:	dt	<=	199	;
						10'd608	:	dt	<=	225	;
						10'd609	:	dt	<=	224	;
						10'd610	:	dt	<=	222	;
						10'd611	:	dt	<=	191	;
						10'd612	:	dt	<=	125	;
						10'd613	:	dt	<=	164	;
						10'd614	:	dt	<=	255	;
						10'd615	:	dt	<=	250	;
						10'd616	:	dt	<=	120	;
						10'd617	:	dt	<=	122	;
						10'd618	:	dt	<=	130	;
						10'd619	:	dt	<=	147	;
						10'd620	:	dt	<=	160	;
						10'd621	:	dt	<=	160	;
						10'd622	:	dt	<=	103	;
						10'd623	:	dt	<=	100	;
						10'd624	:	dt	<=	79	;
						10'd625	:	dt	<=	104	;
						10'd626	:	dt	<=	108	;
						10'd627	:	dt	<=	117	;
						10'd628	:	dt	<=	108	;
						10'd629	:	dt	<=	80	;
						10'd630	:	dt	<=	66	;
						10'd631	:	dt	<=	93	;
						10'd632	:	dt	<=	107	;
						10'd633	:	dt	<=	117	;
						10'd634	:	dt	<=	104	;
						10'd635	:	dt	<=	84	;
						10'd636	:	dt	<=	115	;
						10'd637	:	dt	<=	179	;
						10'd638	:	dt	<=	194	;
						10'd639	:	dt	<=	167	;
						10'd640	:	dt	<=	184	;
						10'd641	:	dt	<=	250	;
						10'd642	:	dt	<=	255	;
						10'd643	:	dt	<=	253	;
						10'd644	:	dt	<=	120	;
						10'd645	:	dt	<=	121	;
						10'd646	:	dt	<=	131	;
						10'd647	:	dt	<=	147	;
						10'd648	:	dt	<=	168	;
						10'd649	:	dt	<=	153	;
						10'd650	:	dt	<=	88	;
						10'd651	:	dt	<=	89	;
						10'd652	:	dt	<=	75	;
						10'd653	:	dt	<=	84	;
						10'd654	:	dt	<=	178	;
						10'd655	:	dt	<=	138	;
						10'd656	:	dt	<=	105	;
						10'd657	:	dt	<=	94	;
						10'd658	:	dt	<=	74	;
						10'd659	:	dt	<=	58	;
						10'd660	:	dt	<=	58	;
						10'd661	:	dt	<=	46	;
						10'd662	:	dt	<=	44	;
						10'd663	:	dt	<=	44	;
						10'd664	:	dt	<=	11	;
						10'd665	:	dt	<=	119	;
						10'd666	:	dt	<=	255	;
						10'd667	:	dt	<=	245	;
						10'd668	:	dt	<=	255	;
						10'd669	:	dt	<=	255	;
						10'd670	:	dt	<=	254	;
						10'd671	:	dt	<=	255	;
						10'd672	:	dt	<=	119	;
						10'd673	:	dt	<=	121	;
						10'd674	:	dt	<=	131	;
						10'd675	:	dt	<=	147	;
						10'd676	:	dt	<=	167	;
						10'd677	:	dt	<=	127	;
						10'd678	:	dt	<=	91	;
						10'd679	:	dt	<=	83	;
						10'd680	:	dt	<=	87	;
						10'd681	:	dt	<=	66	;
						10'd682	:	dt	<=	39	;
						10'd683	:	dt	<=	70	;
						10'd684	:	dt	<=	43	;
						10'd685	:	dt	<=	26	;
						10'd686	:	dt	<=	14	;
						10'd687	:	dt	<=	9	;
						10'd688	:	dt	<=	9	;
						10'd689	:	dt	<=	12	;
						10'd690	:	dt	<=	11	;
						10'd691	:	dt	<=	15	;
						10'd692	:	dt	<=	0	;
						10'd693	:	dt	<=	83	;
						10'd694	:	dt	<=	255	;
						10'd695	:	dt	<=	252	;
						10'd696	:	dt	<=	254	;
						10'd697	:	dt	<=	255	;
						10'd698	:	dt	<=	255	;
						10'd699	:	dt	<=	255	;
						10'd700	:	dt	<=	119	;
						10'd701	:	dt	<=	122	;
						10'd702	:	dt	<=	131	;
						10'd703	:	dt	<=	152	;
						10'd704	:	dt	<=	154	;
						10'd705	:	dt	<=	106	;
						10'd706	:	dt	<=	89	;
						10'd707	:	dt	<=	80	;
						10'd708	:	dt	<=	74	;
						10'd709	:	dt	<=	91	;
						10'd710	:	dt	<=	31	;
						10'd711	:	dt	<=	0	;
						10'd712	:	dt	<=	30	;
						10'd713	:	dt	<=	26	;
						10'd714	:	dt	<=	16	;
						10'd715	:	dt	<=	8	;
						10'd716	:	dt	<=	8	;
						10'd717	:	dt	<=	9	;
						10'd718	:	dt	<=	10	;
						10'd719	:	dt	<=	12	;
						10'd720	:	dt	<=	0	;
						10'd721	:	dt	<=	193	;
						10'd722	:	dt	<=	255	;
						10'd723	:	dt	<=	250	;
						10'd724	:	dt	<=	255	;
						10'd725	:	dt	<=	255	;
						10'd726	:	dt	<=	255	;
						10'd727	:	dt	<=	255	;
						10'd728	:	dt	<=	118	;
						10'd729	:	dt	<=	121	;
						10'd730	:	dt	<=	131	;
						10'd731	:	dt	<=	153	;
						10'd732	:	dt	<=	133	;
						10'd733	:	dt	<=	95	;
						10'd734	:	dt	<=	85	;
						10'd735	:	dt	<=	76	;
						10'd736	:	dt	<=	72	;
						10'd737	:	dt	<=	76	;
						10'd738	:	dt	<=	69	;
						10'd739	:	dt	<=	0	;
						10'd740	:	dt	<=	17	;
						10'd741	:	dt	<=	29	;
						10'd742	:	dt	<=	17	;
						10'd743	:	dt	<=	9	;
						10'd744	:	dt	<=	8	;
						10'd745	:	dt	<=	8	;
						10'd746	:	dt	<=	11	;
						10'd747	:	dt	<=	1	;
						10'd748	:	dt	<=	36	;
						10'd749	:	dt	<=	252	;
						10'd750	:	dt	<=	253	;
						10'd751	:	dt	<=	254	;
						10'd752	:	dt	<=	255	;
						10'd753	:	dt	<=	255	;
						10'd754	:	dt	<=	255	;
						10'd755	:	dt	<=	255	;
						10'd756	:	dt	<=	117	;
						10'd757	:	dt	<=	122	;
						10'd758	:	dt	<=	132	;
						10'd759	:	dt	<=	149	;
						10'd760	:	dt	<=	106	;
						10'd761	:	dt	<=	87	;
						10'd762	:	dt	<=	83	;
						10'd763	:	dt	<=	74	;
						10'd764	:	dt	<=	68	;
						10'd765	:	dt	<=	73	;
						10'd766	:	dt	<=	80	;
						10'd767	:	dt	<=	6	;
						10'd768	:	dt	<=	0	;
						10'd769	:	dt	<=	22	;
						10'd770	:	dt	<=	16	;
						10'd771	:	dt	<=	10	;
						10'd772	:	dt	<=	8	;
						10'd773	:	dt	<=	7	;
						10'd774	:	dt	<=	12	;
						10'd775	:	dt	<=	0	;
						10'd776	:	dt	<=	104	;
						10'd777	:	dt	<=	255	;
						10'd778	:	dt	<=	251	;
						10'd779	:	dt	<=	255	;
						10'd780	:	dt	<=	255	;
						10'd781	:	dt	<=	255	;
						10'd782	:	dt	<=	255	;
						10'd783	:	dt	<=	255	;
					endcase
				end
				5'd17	:	begin
					case (cnt)
						10'd0	:	dt	<=	138	;
						10'd1	:	dt	<=	139	;
						10'd2	:	dt	<=	141	;
						10'd3	:	dt	<=	143	;
						10'd4	:	dt	<=	147	;
						10'd5	:	dt	<=	149	;
						10'd6	:	dt	<=	149	;
						10'd7	:	dt	<=	152	;
						10'd8	:	dt	<=	153	;
						10'd9	:	dt	<=	153	;
						10'd10	:	dt	<=	154	;
						10'd11	:	dt	<=	156	;
						10'd12	:	dt	<=	157	;
						10'd13	:	dt	<=	158	;
						10'd14	:	dt	<=	160	;
						10'd15	:	dt	<=	161	;
						10'd16	:	dt	<=	161	;
						10'd17	:	dt	<=	161	;
						10'd18	:	dt	<=	162	;
						10'd19	:	dt	<=	162	;
						10'd20	:	dt	<=	164	;
						10'd21	:	dt	<=	163	;
						10'd22	:	dt	<=	163	;
						10'd23	:	dt	<=	163	;
						10'd24	:	dt	<=	162	;
						10'd25	:	dt	<=	163	;
						10'd26	:	dt	<=	164	;
						10'd27	:	dt	<=	163	;
						10'd28	:	dt	<=	139	;
						10'd29	:	dt	<=	140	;
						10'd30	:	dt	<=	142	;
						10'd31	:	dt	<=	146	;
						10'd32	:	dt	<=	148	;
						10'd33	:	dt	<=	149	;
						10'd34	:	dt	<=	150	;
						10'd35	:	dt	<=	153	;
						10'd36	:	dt	<=	153	;
						10'd37	:	dt	<=	154	;
						10'd38	:	dt	<=	156	;
						10'd39	:	dt	<=	157	;
						10'd40	:	dt	<=	158	;
						10'd41	:	dt	<=	160	;
						10'd42	:	dt	<=	160	;
						10'd43	:	dt	<=	162	;
						10'd44	:	dt	<=	162	;
						10'd45	:	dt	<=	162	;
						10'd46	:	dt	<=	163	;
						10'd47	:	dt	<=	163	;
						10'd48	:	dt	<=	164	;
						10'd49	:	dt	<=	164	;
						10'd50	:	dt	<=	165	;
						10'd51	:	dt	<=	166	;
						10'd52	:	dt	<=	165	;
						10'd53	:	dt	<=	166	;
						10'd54	:	dt	<=	166	;
						10'd55	:	dt	<=	165	;
						10'd56	:	dt	<=	140	;
						10'd57	:	dt	<=	142	;
						10'd58	:	dt	<=	145	;
						10'd59	:	dt	<=	148	;
						10'd60	:	dt	<=	150	;
						10'd61	:	dt	<=	151	;
						10'd62	:	dt	<=	152	;
						10'd63	:	dt	<=	154	;
						10'd64	:	dt	<=	155	;
						10'd65	:	dt	<=	156	;
						10'd66	:	dt	<=	158	;
						10'd67	:	dt	<=	158	;
						10'd68	:	dt	<=	159	;
						10'd69	:	dt	<=	161	;
						10'd70	:	dt	<=	162	;
						10'd71	:	dt	<=	162	;
						10'd72	:	dt	<=	163	;
						10'd73	:	dt	<=	165	;
						10'd74	:	dt	<=	164	;
						10'd75	:	dt	<=	164	;
						10'd76	:	dt	<=	166	;
						10'd77	:	dt	<=	165	;
						10'd78	:	dt	<=	166	;
						10'd79	:	dt	<=	167	;
						10'd80	:	dt	<=	167	;
						10'd81	:	dt	<=	167	;
						10'd82	:	dt	<=	168	;
						10'd83	:	dt	<=	167	;
						10'd84	:	dt	<=	142	;
						10'd85	:	dt	<=	143	;
						10'd86	:	dt	<=	147	;
						10'd87	:	dt	<=	148	;
						10'd88	:	dt	<=	150	;
						10'd89	:	dt	<=	152	;
						10'd90	:	dt	<=	153	;
						10'd91	:	dt	<=	154	;
						10'd92	:	dt	<=	156	;
						10'd93	:	dt	<=	157	;
						10'd94	:	dt	<=	159	;
						10'd95	:	dt	<=	159	;
						10'd96	:	dt	<=	161	;
						10'd97	:	dt	<=	162	;
						10'd98	:	dt	<=	164	;
						10'd99	:	dt	<=	163	;
						10'd100	:	dt	<=	165	;
						10'd101	:	dt	<=	167	;
						10'd102	:	dt	<=	166	;
						10'd103	:	dt	<=	167	;
						10'd104	:	dt	<=	169	;
						10'd105	:	dt	<=	167	;
						10'd106	:	dt	<=	167	;
						10'd107	:	dt	<=	169	;
						10'd108	:	dt	<=	167	;
						10'd109	:	dt	<=	168	;
						10'd110	:	dt	<=	168	;
						10'd111	:	dt	<=	168	;
						10'd112	:	dt	<=	141	;
						10'd113	:	dt	<=	144	;
						10'd114	:	dt	<=	147	;
						10'd115	:	dt	<=	149	;
						10'd116	:	dt	<=	151	;
						10'd117	:	dt	<=	153	;
						10'd118	:	dt	<=	154	;
						10'd119	:	dt	<=	155	;
						10'd120	:	dt	<=	157	;
						10'd121	:	dt	<=	158	;
						10'd122	:	dt	<=	160	;
						10'd123	:	dt	<=	161	;
						10'd124	:	dt	<=	162	;
						10'd125	:	dt	<=	164	;
						10'd126	:	dt	<=	164	;
						10'd127	:	dt	<=	166	;
						10'd128	:	dt	<=	167	;
						10'd129	:	dt	<=	167	;
						10'd130	:	dt	<=	163	;
						10'd131	:	dt	<=	171	;
						10'd132	:	dt	<=	167	;
						10'd133	:	dt	<=	168	;
						10'd134	:	dt	<=	169	;
						10'd135	:	dt	<=	169	;
						10'd136	:	dt	<=	168	;
						10'd137	:	dt	<=	169	;
						10'd138	:	dt	<=	170	;
						10'd139	:	dt	<=	169	;
						10'd140	:	dt	<=	142	;
						10'd141	:	dt	<=	144	;
						10'd142	:	dt	<=	147	;
						10'd143	:	dt	<=	149	;
						10'd144	:	dt	<=	152	;
						10'd145	:	dt	<=	154	;
						10'd146	:	dt	<=	155	;
						10'd147	:	dt	<=	156	;
						10'd148	:	dt	<=	158	;
						10'd149	:	dt	<=	158	;
						10'd150	:	dt	<=	161	;
						10'd151	:	dt	<=	163	;
						10'd152	:	dt	<=	163	;
						10'd153	:	dt	<=	163	;
						10'd154	:	dt	<=	166	;
						10'd155	:	dt	<=	167	;
						10'd156	:	dt	<=	166	;
						10'd157	:	dt	<=	170	;
						10'd158	:	dt	<=	148	;
						10'd159	:	dt	<=	126	;
						10'd160	:	dt	<=	127	;
						10'd161	:	dt	<=	121	;
						10'd162	:	dt	<=	174	;
						10'd163	:	dt	<=	169	;
						10'd164	:	dt	<=	170	;
						10'd165	:	dt	<=	170	;
						10'd166	:	dt	<=	171	;
						10'd167	:	dt	<=	170	;
						10'd168	:	dt	<=	143	;
						10'd169	:	dt	<=	145	;
						10'd170	:	dt	<=	148	;
						10'd171	:	dt	<=	150	;
						10'd172	:	dt	<=	152	;
						10'd173	:	dt	<=	155	;
						10'd174	:	dt	<=	156	;
						10'd175	:	dt	<=	158	;
						10'd176	:	dt	<=	159	;
						10'd177	:	dt	<=	161	;
						10'd178	:	dt	<=	162	;
						10'd179	:	dt	<=	163	;
						10'd180	:	dt	<=	163	;
						10'd181	:	dt	<=	165	;
						10'd182	:	dt	<=	167	;
						10'd183	:	dt	<=	168	;
						10'd184	:	dt	<=	166	;
						10'd185	:	dt	<=	177	;
						10'd186	:	dt	<=	172	;
						10'd187	:	dt	<=	108	;
						10'd188	:	dt	<=	78	;
						10'd189	:	dt	<=	99	;
						10'd190	:	dt	<=	173	;
						10'd191	:	dt	<=	170	;
						10'd192	:	dt	<=	171	;
						10'd193	:	dt	<=	171	;
						10'd194	:	dt	<=	171	;
						10'd195	:	dt	<=	171	;
						10'd196	:	dt	<=	145	;
						10'd197	:	dt	<=	146	;
						10'd198	:	dt	<=	149	;
						10'd199	:	dt	<=	152	;
						10'd200	:	dt	<=	153	;
						10'd201	:	dt	<=	155	;
						10'd202	:	dt	<=	156	;
						10'd203	:	dt	<=	159	;
						10'd204	:	dt	<=	161	;
						10'd205	:	dt	<=	164	;
						10'd206	:	dt	<=	164	;
						10'd207	:	dt	<=	165	;
						10'd208	:	dt	<=	166	;
						10'd209	:	dt	<=	168	;
						10'd210	:	dt	<=	167	;
						10'd211	:	dt	<=	168	;
						10'd212	:	dt	<=	168	;
						10'd213	:	dt	<=	177	;
						10'd214	:	dt	<=	181	;
						10'd215	:	dt	<=	129	;
						10'd216	:	dt	<=	71	;
						10'd217	:	dt	<=	107	;
						10'd218	:	dt	<=	181	;
						10'd219	:	dt	<=	170	;
						10'd220	:	dt	<=	172	;
						10'd221	:	dt	<=	172	;
						10'd222	:	dt	<=	171	;
						10'd223	:	dt	<=	172	;
						10'd224	:	dt	<=	146	;
						10'd225	:	dt	<=	147	;
						10'd226	:	dt	<=	149	;
						10'd227	:	dt	<=	152	;
						10'd228	:	dt	<=	154	;
						10'd229	:	dt	<=	155	;
						10'd230	:	dt	<=	158	;
						10'd231	:	dt	<=	160	;
						10'd232	:	dt	<=	162	;
						10'd233	:	dt	<=	163	;
						10'd234	:	dt	<=	164	;
						10'd235	:	dt	<=	166	;
						10'd236	:	dt	<=	167	;
						10'd237	:	dt	<=	164	;
						10'd238	:	dt	<=	171	;
						10'd239	:	dt	<=	170	;
						10'd240	:	dt	<=	170	;
						10'd241	:	dt	<=	173	;
						10'd242	:	dt	<=	187	;
						10'd243	:	dt	<=	149	;
						10'd244	:	dt	<=	82	;
						10'd245	:	dt	<=	126	;
						10'd246	:	dt	<=	183	;
						10'd247	:	dt	<=	171	;
						10'd248	:	dt	<=	173	;
						10'd249	:	dt	<=	172	;
						10'd250	:	dt	<=	172	;
						10'd251	:	dt	<=	173	;
						10'd252	:	dt	<=	146	;
						10'd253	:	dt	<=	148	;
						10'd254	:	dt	<=	151	;
						10'd255	:	dt	<=	154	;
						10'd256	:	dt	<=	155	;
						10'd257	:	dt	<=	157	;
						10'd258	:	dt	<=	160	;
						10'd259	:	dt	<=	160	;
						10'd260	:	dt	<=	161	;
						10'd261	:	dt	<=	163	;
						10'd262	:	dt	<=	164	;
						10'd263	:	dt	<=	163	;
						10'd264	:	dt	<=	169	;
						10'd265	:	dt	<=	150	;
						10'd266	:	dt	<=	133	;
						10'd267	:	dt	<=	174	;
						10'd268	:	dt	<=	171	;
						10'd269	:	dt	<=	174	;
						10'd270	:	dt	<=	188	;
						10'd271	:	dt	<=	148	;
						10'd272	:	dt	<=	97	;
						10'd273	:	dt	<=	156	;
						10'd274	:	dt	<=	179	;
						10'd275	:	dt	<=	175	;
						10'd276	:	dt	<=	175	;
						10'd277	:	dt	<=	173	;
						10'd278	:	dt	<=	173	;
						10'd279	:	dt	<=	173	;
						10'd280	:	dt	<=	145	;
						10'd281	:	dt	<=	149	;
						10'd282	:	dt	<=	152	;
						10'd283	:	dt	<=	153	;
						10'd284	:	dt	<=	155	;
						10'd285	:	dt	<=	158	;
						10'd286	:	dt	<=	160	;
						10'd287	:	dt	<=	160	;
						10'd288	:	dt	<=	162	;
						10'd289	:	dt	<=	163	;
						10'd290	:	dt	<=	165	;
						10'd291	:	dt	<=	167	;
						10'd292	:	dt	<=	175	;
						10'd293	:	dt	<=	161	;
						10'd294	:	dt	<=	115	;
						10'd295	:	dt	<=	124	;
						10'd296	:	dt	<=	173	;
						10'd297	:	dt	<=	187	;
						10'd298	:	dt	<=	183	;
						10'd299	:	dt	<=	141	;
						10'd300	:	dt	<=	101	;
						10'd301	:	dt	<=	165	;
						10'd302	:	dt	<=	178	;
						10'd303	:	dt	<=	176	;
						10'd304	:	dt	<=	175	;
						10'd305	:	dt	<=	175	;
						10'd306	:	dt	<=	174	;
						10'd307	:	dt	<=	173	;
						10'd308	:	dt	<=	146	;
						10'd309	:	dt	<=	149	;
						10'd310	:	dt	<=	152	;
						10'd311	:	dt	<=	154	;
						10'd312	:	dt	<=	157	;
						10'd313	:	dt	<=	158	;
						10'd314	:	dt	<=	161	;
						10'd315	:	dt	<=	161	;
						10'd316	:	dt	<=	162	;
						10'd317	:	dt	<=	167	;
						10'd318	:	dt	<=	156	;
						10'd319	:	dt	<=	136	;
						10'd320	:	dt	<=	170	;
						10'd321	:	dt	<=	177	;
						10'd322	:	dt	<=	162	;
						10'd323	:	dt	<=	143	;
						10'd324	:	dt	<=	120	;
						10'd325	:	dt	<=	151	;
						10'd326	:	dt	<=	175	;
						10'd327	:	dt	<=	144	;
						10'd328	:	dt	<=	99	;
						10'd329	:	dt	<=	164	;
						10'd330	:	dt	<=	180	;
						10'd331	:	dt	<=	176	;
						10'd332	:	dt	<=	176	;
						10'd333	:	dt	<=	176	;
						10'd334	:	dt	<=	175	;
						10'd335	:	dt	<=	175	;
						10'd336	:	dt	<=	147	;
						10'd337	:	dt	<=	149	;
						10'd338	:	dt	<=	153	;
						10'd339	:	dt	<=	155	;
						10'd340	:	dt	<=	157	;
						10'd341	:	dt	<=	160	;
						10'd342	:	dt	<=	162	;
						10'd343	:	dt	<=	161	;
						10'd344	:	dt	<=	166	;
						10'd345	:	dt	<=	191	;
						10'd346	:	dt	<=	156	;
						10'd347	:	dt	<=	107	;
						10'd348	:	dt	<=	148	;
						10'd349	:	dt	<=	175	;
						10'd350	:	dt	<=	190	;
						10'd351	:	dt	<=	177	;
						10'd352	:	dt	<=	127	;
						10'd353	:	dt	<=	84	;
						10'd354	:	dt	<=	138	;
						10'd355	:	dt	<=	136	;
						10'd356	:	dt	<=	101	;
						10'd357	:	dt	<=	163	;
						10'd358	:	dt	<=	181	;
						10'd359	:	dt	<=	177	;
						10'd360	:	dt	<=	176	;
						10'd361	:	dt	<=	175	;
						10'd362	:	dt	<=	176	;
						10'd363	:	dt	<=	176	;
						10'd364	:	dt	<=	147	;
						10'd365	:	dt	<=	151	;
						10'd366	:	dt	<=	154	;
						10'd367	:	dt	<=	156	;
						10'd368	:	dt	<=	158	;
						10'd369	:	dt	<=	161	;
						10'd370	:	dt	<=	164	;
						10'd371	:	dt	<=	160	;
						10'd372	:	dt	<=	176	;
						10'd373	:	dt	<=	162	;
						10'd374	:	dt	<=	166	;
						10'd375	:	dt	<=	138	;
						10'd376	:	dt	<=	137	;
						10'd377	:	dt	<=	123	;
						10'd378	:	dt	<=	161	;
						10'd379	:	dt	<=	192	;
						10'd380	:	dt	<=	159	;
						10'd381	:	dt	<=	94	;
						10'd382	:	dt	<=	99	;
						10'd383	:	dt	<=	120	;
						10'd384	:	dt	<=	95	;
						10'd385	:	dt	<=	161	;
						10'd386	:	dt	<=	181	;
						10'd387	:	dt	<=	177	;
						10'd388	:	dt	<=	176	;
						10'd389	:	dt	<=	176	;
						10'd390	:	dt	<=	177	;
						10'd391	:	dt	<=	177	;
						10'd392	:	dt	<=	148	;
						10'd393	:	dt	<=	151	;
						10'd394	:	dt	<=	155	;
						10'd395	:	dt	<=	157	;
						10'd396	:	dt	<=	159	;
						10'd397	:	dt	<=	160	;
						10'd398	:	dt	<=	163	;
						10'd399	:	dt	<=	160	;
						10'd400	:	dt	<=	185	;
						10'd401	:	dt	<=	152	;
						10'd402	:	dt	<=	123	;
						10'd403	:	dt	<=	127	;
						10'd404	:	dt	<=	96	;
						10'd405	:	dt	<=	63	;
						10'd406	:	dt	<=	104	;
						10'd407	:	dt	<=	207	;
						10'd408	:	dt	<=	176	;
						10'd409	:	dt	<=	117	;
						10'd410	:	dt	<=	82	;
						10'd411	:	dt	<=	97	;
						10'd412	:	dt	<=	85	;
						10'd413	:	dt	<=	161	;
						10'd414	:	dt	<=	183	;
						10'd415	:	dt	<=	178	;
						10'd416	:	dt	<=	177	;
						10'd417	:	dt	<=	177	;
						10'd418	:	dt	<=	177	;
						10'd419	:	dt	<=	177	;
						10'd420	:	dt	<=	150	;
						10'd421	:	dt	<=	152	;
						10'd422	:	dt	<=	154	;
						10'd423	:	dt	<=	157	;
						10'd424	:	dt	<=	159	;
						10'd425	:	dt	<=	161	;
						10'd426	:	dt	<=	164	;
						10'd427	:	dt	<=	165	;
						10'd428	:	dt	<=	181	;
						10'd429	:	dt	<=	142	;
						10'd430	:	dt	<=	109	;
						10'd431	:	dt	<=	126	;
						10'd432	:	dt	<=	103	;
						10'd433	:	dt	<=	90	;
						10'd434	:	dt	<=	104	;
						10'd435	:	dt	<=	203	;
						10'd436	:	dt	<=	190	;
						10'd437	:	dt	<=	140	;
						10'd438	:	dt	<=	83	;
						10'd439	:	dt	<=	87	;
						10'd440	:	dt	<=	80	;
						10'd441	:	dt	<=	157	;
						10'd442	:	dt	<=	183	;
						10'd443	:	dt	<=	178	;
						10'd444	:	dt	<=	179	;
						10'd445	:	dt	<=	178	;
						10'd446	:	dt	<=	177	;
						10'd447	:	dt	<=	178	;
						10'd448	:	dt	<=	149	;
						10'd449	:	dt	<=	152	;
						10'd450	:	dt	<=	155	;
						10'd451	:	dt	<=	158	;
						10'd452	:	dt	<=	160	;
						10'd453	:	dt	<=	163	;
						10'd454	:	dt	<=	163	;
						10'd455	:	dt	<=	171	;
						10'd456	:	dt	<=	186	;
						10'd457	:	dt	<=	160	;
						10'd458	:	dt	<=	144	;
						10'd459	:	dt	<=	133	;
						10'd460	:	dt	<=	112	;
						10'd461	:	dt	<=	134	;
						10'd462	:	dt	<=	120	;
						10'd463	:	dt	<=	192	;
						10'd464	:	dt	<=	195	;
						10'd465	:	dt	<=	150	;
						10'd466	:	dt	<=	97	;
						10'd467	:	dt	<=	83	;
						10'd468	:	dt	<=	81	;
						10'd469	:	dt	<=	152	;
						10'd470	:	dt	<=	185	;
						10'd471	:	dt	<=	178	;
						10'd472	:	dt	<=	179	;
						10'd473	:	dt	<=	179	;
						10'd474	:	dt	<=	178	;
						10'd475	:	dt	<=	178	;
						10'd476	:	dt	<=	150	;
						10'd477	:	dt	<=	152	;
						10'd478	:	dt	<=	155	;
						10'd479	:	dt	<=	159	;
						10'd480	:	dt	<=	160	;
						10'd481	:	dt	<=	163	;
						10'd482	:	dt	<=	161	;
						10'd483	:	dt	<=	181	;
						10'd484	:	dt	<=	178	;
						10'd485	:	dt	<=	141	;
						10'd486	:	dt	<=	135	;
						10'd487	:	dt	<=	128	;
						10'd488	:	dt	<=	124	;
						10'd489	:	dt	<=	144	;
						10'd490	:	dt	<=	169	;
						10'd491	:	dt	<=	192	;
						10'd492	:	dt	<=	176	;
						10'd493	:	dt	<=	157	;
						10'd494	:	dt	<=	107	;
						10'd495	:	dt	<=	78	;
						10'd496	:	dt	<=	77	;
						10'd497	:	dt	<=	154	;
						10'd498	:	dt	<=	186	;
						10'd499	:	dt	<=	178	;
						10'd500	:	dt	<=	181	;
						10'd501	:	dt	<=	181	;
						10'd502	:	dt	<=	179	;
						10'd503	:	dt	<=	179	;
						10'd504	:	dt	<=	151	;
						10'd505	:	dt	<=	153	;
						10'd506	:	dt	<=	156	;
						10'd507	:	dt	<=	158	;
						10'd508	:	dt	<=	162	;
						10'd509	:	dt	<=	165	;
						10'd510	:	dt	<=	163	;
						10'd511	:	dt	<=	189	;
						10'd512	:	dt	<=	166	;
						10'd513	:	dt	<=	138	;
						10'd514	:	dt	<=	129	;
						10'd515	:	dt	<=	129	;
						10'd516	:	dt	<=	137	;
						10'd517	:	dt	<=	157	;
						10'd518	:	dt	<=	214	;
						10'd519	:	dt	<=	190	;
						10'd520	:	dt	<=	157	;
						10'd521	:	dt	<=	146	;
						10'd522	:	dt	<=	104	;
						10'd523	:	dt	<=	74	;
						10'd524	:	dt	<=	70	;
						10'd525	:	dt	<=	156	;
						10'd526	:	dt	<=	187	;
						10'd527	:	dt	<=	180	;
						10'd528	:	dt	<=	181	;
						10'd529	:	dt	<=	181	;
						10'd530	:	dt	<=	180	;
						10'd531	:	dt	<=	180	;
						10'd532	:	dt	<=	152	;
						10'd533	:	dt	<=	154	;
						10'd534	:	dt	<=	155	;
						10'd535	:	dt	<=	159	;
						10'd536	:	dt	<=	162	;
						10'd537	:	dt	<=	164	;
						10'd538	:	dt	<=	163	;
						10'd539	:	dt	<=	195	;
						10'd540	:	dt	<=	169	;
						10'd541	:	dt	<=	146	;
						10'd542	:	dt	<=	131	;
						10'd543	:	dt	<=	132	;
						10'd544	:	dt	<=	140	;
						10'd545	:	dt	<=	196	;
						10'd546	:	dt	<=	206	;
						10'd547	:	dt	<=	187	;
						10'd548	:	dt	<=	155	;
						10'd549	:	dt	<=	135	;
						10'd550	:	dt	<=	99	;
						10'd551	:	dt	<=	73	;
						10'd552	:	dt	<=	71	;
						10'd553	:	dt	<=	166	;
						10'd554	:	dt	<=	185	;
						10'd555	:	dt	<=	182	;
						10'd556	:	dt	<=	181	;
						10'd557	:	dt	<=	181	;
						10'd558	:	dt	<=	181	;
						10'd559	:	dt	<=	181	;
						10'd560	:	dt	<=	151	;
						10'd561	:	dt	<=	154	;
						10'd562	:	dt	<=	156	;
						10'd563	:	dt	<=	160	;
						10'd564	:	dt	<=	161	;
						10'd565	:	dt	<=	163	;
						10'd566	:	dt	<=	168	;
						10'd567	:	dt	<=	199	;
						10'd568	:	dt	<=	171	;
						10'd569	:	dt	<=	156	;
						10'd570	:	dt	<=	133	;
						10'd571	:	dt	<=	132	;
						10'd572	:	dt	<=	166	;
						10'd573	:	dt	<=	212	;
						10'd574	:	dt	<=	192	;
						10'd575	:	dt	<=	180	;
						10'd576	:	dt	<=	146	;
						10'd577	:	dt	<=	128	;
						10'd578	:	dt	<=	94	;
						10'd579	:	dt	<=	70	;
						10'd580	:	dt	<=	89	;
						10'd581	:	dt	<=	185	;
						10'd582	:	dt	<=	181	;
						10'd583	:	dt	<=	181	;
						10'd584	:	dt	<=	180	;
						10'd585	:	dt	<=	181	;
						10'd586	:	dt	<=	181	;
						10'd587	:	dt	<=	181	;
						10'd588	:	dt	<=	151	;
						10'd589	:	dt	<=	153	;
						10'd590	:	dt	<=	158	;
						10'd591	:	dt	<=	161	;
						10'd592	:	dt	<=	163	;
						10'd593	:	dt	<=	161	;
						10'd594	:	dt	<=	174	;
						10'd595	:	dt	<=	201	;
						10'd596	:	dt	<=	172	;
						10'd597	:	dt	<=	163	;
						10'd598	:	dt	<=	147	;
						10'd599	:	dt	<=	133	;
						10'd600	:	dt	<=	186	;
						10'd601	:	dt	<=	209	;
						10'd602	:	dt	<=	187	;
						10'd603	:	dt	<=	178	;
						10'd604	:	dt	<=	138	;
						10'd605	:	dt	<=	116	;
						10'd606	:	dt	<=	91	;
						10'd607	:	dt	<=	64	;
						10'd608	:	dt	<=	127	;
						10'd609	:	dt	<=	191	;
						10'd610	:	dt	<=	180	;
						10'd611	:	dt	<=	182	;
						10'd612	:	dt	<=	181	;
						10'd613	:	dt	<=	181	;
						10'd614	:	dt	<=	179	;
						10'd615	:	dt	<=	179	;
						10'd616	:	dt	<=	151	;
						10'd617	:	dt	<=	154	;
						10'd618	:	dt	<=	157	;
						10'd619	:	dt	<=	161	;
						10'd620	:	dt	<=	166	;
						10'd621	:	dt	<=	163	;
						10'd622	:	dt	<=	179	;
						10'd623	:	dt	<=	206	;
						10'd624	:	dt	<=	176	;
						10'd625	:	dt	<=	172	;
						10'd626	:	dt	<=	163	;
						10'd627	:	dt	<=	142	;
						10'd628	:	dt	<=	189	;
						10'd629	:	dt	<=	197	;
						10'd630	:	dt	<=	180	;
						10'd631	:	dt	<=	172	;
						10'd632	:	dt	<=	141	;
						10'd633	:	dt	<=	105	;
						10'd634	:	dt	<=	84	;
						10'd635	:	dt	<=	73	;
						10'd636	:	dt	<=	169	;
						10'd637	:	dt	<=	185	;
						10'd638	:	dt	<=	181	;
						10'd639	:	dt	<=	183	;
						10'd640	:	dt	<=	183	;
						10'd641	:	dt	<=	183	;
						10'd642	:	dt	<=	181	;
						10'd643	:	dt	<=	181	;
						10'd644	:	dt	<=	152	;
						10'd645	:	dt	<=	155	;
						10'd646	:	dt	<=	159	;
						10'd647	:	dt	<=	162	;
						10'd648	:	dt	<=	165	;
						10'd649	:	dt	<=	163	;
						10'd650	:	dt	<=	176	;
						10'd651	:	dt	<=	210	;
						10'd652	:	dt	<=	183	;
						10'd653	:	dt	<=	177	;
						10'd654	:	dt	<=	170	;
						10'd655	:	dt	<=	152	;
						10'd656	:	dt	<=	175	;
						10'd657	:	dt	<=	190	;
						10'd658	:	dt	<=	177	;
						10'd659	:	dt	<=	165	;
						10'd660	:	dt	<=	135	;
						10'd661	:	dt	<=	102	;
						10'd662	:	dt	<=	72	;
						10'd663	:	dt	<=	111	;
						10'd664	:	dt	<=	192	;
						10'd665	:	dt	<=	181	;
						10'd666	:	dt	<=	182	;
						10'd667	:	dt	<=	182	;
						10'd668	:	dt	<=	184	;
						10'd669	:	dt	<=	184	;
						10'd670	:	dt	<=	182	;
						10'd671	:	dt	<=	181	;
						10'd672	:	dt	<=	152	;
						10'd673	:	dt	<=	155	;
						10'd674	:	dt	<=	159	;
						10'd675	:	dt	<=	163	;
						10'd676	:	dt	<=	165	;
						10'd677	:	dt	<=	165	;
						10'd678	:	dt	<=	171	;
						10'd679	:	dt	<=	207	;
						10'd680	:	dt	<=	191	;
						10'd681	:	dt	<=	173	;
						10'd682	:	dt	<=	163	;
						10'd683	:	dt	<=	161	;
						10'd684	:	dt	<=	165	;
						10'd685	:	dt	<=	180	;
						10'd686	:	dt	<=	171	;
						10'd687	:	dt	<=	174	;
						10'd688	:	dt	<=	131	;
						10'd689	:	dt	<=	97	;
						10'd690	:	dt	<=	69	;
						10'd691	:	dt	<=	142	;
						10'd692	:	dt	<=	191	;
						10'd693	:	dt	<=	180	;
						10'd694	:	dt	<=	181	;
						10'd695	:	dt	<=	183	;
						10'd696	:	dt	<=	183	;
						10'd697	:	dt	<=	182	;
						10'd698	:	dt	<=	182	;
						10'd699	:	dt	<=	182	;
						10'd700	:	dt	<=	153	;
						10'd701	:	dt	<=	155	;
						10'd702	:	dt	<=	160	;
						10'd703	:	dt	<=	163	;
						10'd704	:	dt	<=	165	;
						10'd705	:	dt	<=	168	;
						10'd706	:	dt	<=	167	;
						10'd707	:	dt	<=	202	;
						10'd708	:	dt	<=	186	;
						10'd709	:	dt	<=	172	;
						10'd710	:	dt	<=	157	;
						10'd711	:	dt	<=	159	;
						10'd712	:	dt	<=	168	;
						10'd713	:	dt	<=	169	;
						10'd714	:	dt	<=	170	;
						10'd715	:	dt	<=	175	;
						10'd716	:	dt	<=	132	;
						10'd717	:	dt	<=	95	;
						10'd718	:	dt	<=	73	;
						10'd719	:	dt	<=	161	;
						10'd720	:	dt	<=	189	;
						10'd721	:	dt	<=	183	;
						10'd722	:	dt	<=	184	;
						10'd723	:	dt	<=	184	;
						10'd724	:	dt	<=	184	;
						10'd725	:	dt	<=	183	;
						10'd726	:	dt	<=	183	;
						10'd727	:	dt	<=	184	;
						10'd728	:	dt	<=	153	;
						10'd729	:	dt	<=	156	;
						10'd730	:	dt	<=	159	;
						10'd731	:	dt	<=	161	;
						10'd732	:	dt	<=	164	;
						10'd733	:	dt	<=	166	;
						10'd734	:	dt	<=	170	;
						10'd735	:	dt	<=	201	;
						10'd736	:	dt	<=	184	;
						10'd737	:	dt	<=	173	;
						10'd738	:	dt	<=	158	;
						10'd739	:	dt	<=	158	;
						10'd740	:	dt	<=	168	;
						10'd741	:	dt	<=	166	;
						10'd742	:	dt	<=	170	;
						10'd743	:	dt	<=	166	;
						10'd744	:	dt	<=	123	;
						10'd745	:	dt	<=	91	;
						10'd746	:	dt	<=	94	;
						10'd747	:	dt	<=	184	;
						10'd748	:	dt	<=	185	;
						10'd749	:	dt	<=	184	;
						10'd750	:	dt	<=	185	;
						10'd751	:	dt	<=	185	;
						10'd752	:	dt	<=	184	;
						10'd753	:	dt	<=	184	;
						10'd754	:	dt	<=	184	;
						10'd755	:	dt	<=	183	;
						10'd756	:	dt	<=	152	;
						10'd757	:	dt	<=	154	;
						10'd758	:	dt	<=	157	;
						10'd759	:	dt	<=	161	;
						10'd760	:	dt	<=	165	;
						10'd761	:	dt	<=	165	;
						10'd762	:	dt	<=	174	;
						10'd763	:	dt	<=	203	;
						10'd764	:	dt	<=	194	;
						10'd765	:	dt	<=	175	;
						10'd766	:	dt	<=	164	;
						10'd767	:	dt	<=	167	;
						10'd768	:	dt	<=	174	;
						10'd769	:	dt	<=	160	;
						10'd770	:	dt	<=	166	;
						10'd771	:	dt	<=	153	;
						10'd772	:	dt	<=	112	;
						10'd773	:	dt	<=	80	;
						10'd774	:	dt	<=	136	;
						10'd775	:	dt	<=	193	;
						10'd776	:	dt	<=	183	;
						10'd777	:	dt	<=	184	;
						10'd778	:	dt	<=	184	;
						10'd779	:	dt	<=	184	;
						10'd780	:	dt	<=	184	;
						10'd781	:	dt	<=	185	;
						10'd782	:	dt	<=	185	;
						10'd783	:	dt	<=	183	;
					endcase
				end
				5'd18	:	begin
					case (cnt)
						10'd0	:	dt	<=	198	;
						10'd1	:	dt	<=	202	;
						10'd2	:	dt	<=	204	;
						10'd3	:	dt	<=	204	;
						10'd4	:	dt	<=	206	;
						10'd5	:	dt	<=	208	;
						10'd6	:	dt	<=	210	;
						10'd7	:	dt	<=	212	;
						10'd8	:	dt	<=	212	;
						10'd9	:	dt	<=	213	;
						10'd10	:	dt	<=	214	;
						10'd11	:	dt	<=	217	;
						10'd12	:	dt	<=	218	;
						10'd13	:	dt	<=	218	;
						10'd14	:	dt	<=	219	;
						10'd15	:	dt	<=	221	;
						10'd16	:	dt	<=	221	;
						10'd17	:	dt	<=	222	;
						10'd18	:	dt	<=	222	;
						10'd19	:	dt	<=	224	;
						10'd20	:	dt	<=	224	;
						10'd21	:	dt	<=	224	;
						10'd22	:	dt	<=	225	;
						10'd23	:	dt	<=	223	;
						10'd24	:	dt	<=	222	;
						10'd25	:	dt	<=	223	;
						10'd26	:	dt	<=	223	;
						10'd27	:	dt	<=	223	;
						10'd28	:	dt	<=	200	;
						10'd29	:	dt	<=	202	;
						10'd30	:	dt	<=	205	;
						10'd31	:	dt	<=	206	;
						10'd32	:	dt	<=	207	;
						10'd33	:	dt	<=	209	;
						10'd34	:	dt	<=	211	;
						10'd35	:	dt	<=	212	;
						10'd36	:	dt	<=	214	;
						10'd37	:	dt	<=	215	;
						10'd38	:	dt	<=	216	;
						10'd39	:	dt	<=	217	;
						10'd40	:	dt	<=	218	;
						10'd41	:	dt	<=	219	;
						10'd42	:	dt	<=	220	;
						10'd43	:	dt	<=	222	;
						10'd44	:	dt	<=	223	;
						10'd45	:	dt	<=	222	;
						10'd46	:	dt	<=	222	;
						10'd47	:	dt	<=	223	;
						10'd48	:	dt	<=	225	;
						10'd49	:	dt	<=	225	;
						10'd50	:	dt	<=	227	;
						10'd51	:	dt	<=	226	;
						10'd52	:	dt	<=	225	;
						10'd53	:	dt	<=	225	;
						10'd54	:	dt	<=	223	;
						10'd55	:	dt	<=	224	;
						10'd56	:	dt	<=	201	;
						10'd57	:	dt	<=	203	;
						10'd58	:	dt	<=	205	;
						10'd59	:	dt	<=	208	;
						10'd60	:	dt	<=	210	;
						10'd61	:	dt	<=	211	;
						10'd62	:	dt	<=	211	;
						10'd63	:	dt	<=	214	;
						10'd64	:	dt	<=	214	;
						10'd65	:	dt	<=	215	;
						10'd66	:	dt	<=	217	;
						10'd67	:	dt	<=	217	;
						10'd68	:	dt	<=	217	;
						10'd69	:	dt	<=	219	;
						10'd70	:	dt	<=	220	;
						10'd71	:	dt	<=	225	;
						10'd72	:	dt	<=	227	;
						10'd73	:	dt	<=	222	;
						10'd74	:	dt	<=	222	;
						10'd75	:	dt	<=	224	;
						10'd76	:	dt	<=	223	;
						10'd77	:	dt	<=	224	;
						10'd78	:	dt	<=	227	;
						10'd79	:	dt	<=	227	;
						10'd80	:	dt	<=	227	;
						10'd81	:	dt	<=	225	;
						10'd82	:	dt	<=	224	;
						10'd83	:	dt	<=	224	;
						10'd84	:	dt	<=	202	;
						10'd85	:	dt	<=	203	;
						10'd86	:	dt	<=	208	;
						10'd87	:	dt	<=	209	;
						10'd88	:	dt	<=	210	;
						10'd89	:	dt	<=	212	;
						10'd90	:	dt	<=	211	;
						10'd91	:	dt	<=	214	;
						10'd92	:	dt	<=	216	;
						10'd93	:	dt	<=	216	;
						10'd94	:	dt	<=	218	;
						10'd95	:	dt	<=	218	;
						10'd96	:	dt	<=	220	;
						10'd97	:	dt	<=	220	;
						10'd98	:	dt	<=	222	;
						10'd99	:	dt	<=	210	;
						10'd100	:	dt	<=	204	;
						10'd101	:	dt	<=	229	;
						10'd102	:	dt	<=	223	;
						10'd103	:	dt	<=	227	;
						10'd104	:	dt	<=	226	;
						10'd105	:	dt	<=	225	;
						10'd106	:	dt	<=	228	;
						10'd107	:	dt	<=	227	;
						10'd108	:	dt	<=	227	;
						10'd109	:	dt	<=	227	;
						10'd110	:	dt	<=	227	;
						10'd111	:	dt	<=	226	;
						10'd112	:	dt	<=	202	;
						10'd113	:	dt	<=	204	;
						10'd114	:	dt	<=	210	;
						10'd115	:	dt	<=	208	;
						10'd116	:	dt	<=	209	;
						10'd117	:	dt	<=	211	;
						10'd118	:	dt	<=	213	;
						10'd119	:	dt	<=	214	;
						10'd120	:	dt	<=	216	;
						10'd121	:	dt	<=	218	;
						10'd122	:	dt	<=	219	;
						10'd123	:	dt	<=	221	;
						10'd124	:	dt	<=	225	;
						10'd125	:	dt	<=	221	;
						10'd126	:	dt	<=	234	;
						10'd127	:	dt	<=	207	;
						10'd128	:	dt	<=	153	;
						10'd129	:	dt	<=	192	;
						10'd130	:	dt	<=	231	;
						10'd131	:	dt	<=	225	;
						10'd132	:	dt	<=	226	;
						10'd133	:	dt	<=	230	;
						10'd134	:	dt	<=	226	;
						10'd135	:	dt	<=	225	;
						10'd136	:	dt	<=	227	;
						10'd137	:	dt	<=	227	;
						10'd138	:	dt	<=	228	;
						10'd139	:	dt	<=	228	;
						10'd140	:	dt	<=	202	;
						10'd141	:	dt	<=	205	;
						10'd142	:	dt	<=	209	;
						10'd143	:	dt	<=	209	;
						10'd144	:	dt	<=	210	;
						10'd145	:	dt	<=	211	;
						10'd146	:	dt	<=	214	;
						10'd147	:	dt	<=	215	;
						10'd148	:	dt	<=	215	;
						10'd149	:	dt	<=	219	;
						10'd150	:	dt	<=	221	;
						10'd151	:	dt	<=	213	;
						10'd152	:	dt	<=	196	;
						10'd153	:	dt	<=	219	;
						10'd154	:	dt	<=	226	;
						10'd155	:	dt	<=	220	;
						10'd156	:	dt	<=	158	;
						10'd157	:	dt	<=	110	;
						10'd158	:	dt	<=	204	;
						10'd159	:	dt	<=	230	;
						10'd160	:	dt	<=	205	;
						10'd161	:	dt	<=	193	;
						10'd162	:	dt	<=	221	;
						10'd163	:	dt	<=	230	;
						10'd164	:	dt	<=	228	;
						10'd165	:	dt	<=	229	;
						10'd166	:	dt	<=	227	;
						10'd167	:	dt	<=	227	;
						10'd168	:	dt	<=	202	;
						10'd169	:	dt	<=	203	;
						10'd170	:	dt	<=	207	;
						10'd171	:	dt	<=	209	;
						10'd172	:	dt	<=	211	;
						10'd173	:	dt	<=	211	;
						10'd174	:	dt	<=	216	;
						10'd175	:	dt	<=	218	;
						10'd176	:	dt	<=	218	;
						10'd177	:	dt	<=	222	;
						10'd178	:	dt	<=	237	;
						10'd179	:	dt	<=	215	;
						10'd180	:	dt	<=	170	;
						10'd181	:	dt	<=	173	;
						10'd182	:	dt	<=	232	;
						10'd183	:	dt	<=	202	;
						10'd184	:	dt	<=	175	;
						10'd185	:	dt	<=	125	;
						10'd186	:	dt	<=	141	;
						10'd187	:	dt	<=	186	;
						10'd188	:	dt	<=	177	;
						10'd189	:	dt	<=	158	;
						10'd190	:	dt	<=	161	;
						10'd191	:	dt	<=	237	;
						10'd192	:	dt	<=	228	;
						10'd193	:	dt	<=	229	;
						10'd194	:	dt	<=	228	;
						10'd195	:	dt	<=	228	;
						10'd196	:	dt	<=	202	;
						10'd197	:	dt	<=	204	;
						10'd198	:	dt	<=	208	;
						10'd199	:	dt	<=	210	;
						10'd200	:	dt	<=	210	;
						10'd201	:	dt	<=	212	;
						10'd202	:	dt	<=	214	;
						10'd203	:	dt	<=	213	;
						10'd204	:	dt	<=	206	;
						10'd205	:	dt	<=	238	;
						10'd206	:	dt	<=	239	;
						10'd207	:	dt	<=	215	;
						10'd208	:	dt	<=	178	;
						10'd209	:	dt	<=	153	;
						10'd210	:	dt	<=	249	;
						10'd211	:	dt	<=	221	;
						10'd212	:	dt	<=	205	;
						10'd213	:	dt	<=	167	;
						10'd214	:	dt	<=	126	;
						10'd215	:	dt	<=	133	;
						10'd216	:	dt	<=	161	;
						10'd217	:	dt	<=	155	;
						10'd218	:	dt	<=	115	;
						10'd219	:	dt	<=	215	;
						10'd220	:	dt	<=	233	;
						10'd221	:	dt	<=	229	;
						10'd222	:	dt	<=	229	;
						10'd223	:	dt	<=	228	;
						10'd224	:	dt	<=	204	;
						10'd225	:	dt	<=	206	;
						10'd226	:	dt	<=	209	;
						10'd227	:	dt	<=	211	;
						10'd228	:	dt	<=	211	;
						10'd229	:	dt	<=	210	;
						10'd230	:	dt	<=	229	;
						10'd231	:	dt	<=	218	;
						10'd232	:	dt	<=	167	;
						10'd233	:	dt	<=	214	;
						10'd234	:	dt	<=	242	;
						10'd235	:	dt	<=	208	;
						10'd236	:	dt	<=	174	;
						10'd237	:	dt	<=	173	;
						10'd238	:	dt	<=	247	;
						10'd239	:	dt	<=	246	;
						10'd240	:	dt	<=	226	;
						10'd241	:	dt	<=	177	;
						10'd242	:	dt	<=	132	;
						10'd243	:	dt	<=	116	;
						10'd244	:	dt	<=	143	;
						10'd245	:	dt	<=	144	;
						10'd246	:	dt	<=	105	;
						10'd247	:	dt	<=	183	;
						10'd248	:	dt	<=	241	;
						10'd249	:	dt	<=	228	;
						10'd250	:	dt	<=	230	;
						10'd251	:	dt	<=	229	;
						10'd252	:	dt	<=	205	;
						10'd253	:	dt	<=	206	;
						10'd254	:	dt	<=	209	;
						10'd255	:	dt	<=	212	;
						10'd256	:	dt	<=	208	;
						10'd257	:	dt	<=	226	;
						10'd258	:	dt	<=	251	;
						10'd259	:	dt	<=	218	;
						10'd260	:	dt	<=	163	;
						10'd261	:	dt	<=	197	;
						10'd262	:	dt	<=	243	;
						10'd263	:	dt	<=	208	;
						10'd264	:	dt	<=	163	;
						10'd265	:	dt	<=	193	;
						10'd266	:	dt	<=	236	;
						10'd267	:	dt	<=	239	;
						10'd268	:	dt	<=	223	;
						10'd269	:	dt	<=	177	;
						10'd270	:	dt	<=	127	;
						10'd271	:	dt	<=	102	;
						10'd272	:	dt	<=	122	;
						10'd273	:	dt	<=	134	;
						10'd274	:	dt	<=	100	;
						10'd275	:	dt	<=	184	;
						10'd276	:	dt	<=	242	;
						10'd277	:	dt	<=	228	;
						10'd278	:	dt	<=	231	;
						10'd279	:	dt	<=	230	;
						10'd280	:	dt	<=	206	;
						10'd281	:	dt	<=	208	;
						10'd282	:	dt	<=	209	;
						10'd283	:	dt	<=	211	;
						10'd284	:	dt	<=	209	;
						10'd285	:	dt	<=	235	;
						10'd286	:	dt	<=	254	;
						10'd287	:	dt	<=	219	;
						10'd288	:	dt	<=	164	;
						10'd289	:	dt	<=	184	;
						10'd290	:	dt	<=	243	;
						10'd291	:	dt	<=	212	;
						10'd292	:	dt	<=	152	;
						10'd293	:	dt	<=	208	;
						10'd294	:	dt	<=	236	;
						10'd295	:	dt	<=	237	;
						10'd296	:	dt	<=	219	;
						10'd297	:	dt	<=	174	;
						10'd298	:	dt	<=	126	;
						10'd299	:	dt	<=	92	;
						10'd300	:	dt	<=	108	;
						10'd301	:	dt	<=	119	;
						10'd302	:	dt	<=	100	;
						10'd303	:	dt	<=	203	;
						10'd304	:	dt	<=	239	;
						10'd305	:	dt	<=	229	;
						10'd306	:	dt	<=	231	;
						10'd307	:	dt	<=	231	;
						10'd308	:	dt	<=	207	;
						10'd309	:	dt	<=	209	;
						10'd310	:	dt	<=	210	;
						10'd311	:	dt	<=	211	;
						10'd312	:	dt	<=	213	;
						10'd313	:	dt	<=	225	;
						10'd314	:	dt	<=	243	;
						10'd315	:	dt	<=	222	;
						10'd316	:	dt	<=	168	;
						10'd317	:	dt	<=	171	;
						10'd318	:	dt	<=	242	;
						10'd319	:	dt	<=	209	;
						10'd320	:	dt	<=	138	;
						10'd321	:	dt	<=	171	;
						10'd322	:	dt	<=	220	;
						10'd323	:	dt	<=	246	;
						10'd324	:	dt	<=	214	;
						10'd325	:	dt	<=	167	;
						10'd326	:	dt	<=	121	;
						10'd327	:	dt	<=	93	;
						10'd328	:	dt	<=	99	;
						10'd329	:	dt	<=	102	;
						10'd330	:	dt	<=	116	;
						10'd331	:	dt	<=	223	;
						10'd332	:	dt	<=	235	;
						10'd333	:	dt	<=	230	;
						10'd334	:	dt	<=	232	;
						10'd335	:	dt	<=	231	;
						10'd336	:	dt	<=	207	;
						10'd337	:	dt	<=	209	;
						10'd338	:	dt	<=	212	;
						10'd339	:	dt	<=	208	;
						10'd340	:	dt	<=	220	;
						10'd341	:	dt	<=	239	;
						10'd342	:	dt	<=	221	;
						10'd343	:	dt	<=	219	;
						10'd344	:	dt	<=	179	;
						10'd345	:	dt	<=	152	;
						10'd346	:	dt	<=	219	;
						10'd347	:	dt	<=	195	;
						10'd348	:	dt	<=	137	;
						10'd349	:	dt	<=	94	;
						10'd350	:	dt	<=	186	;
						10'd351	:	dt	<=	253	;
						10'd352	:	dt	<=	205	;
						10'd353	:	dt	<=	161	;
						10'd354	:	dt	<=	115	;
						10'd355	:	dt	<=	96	;
						10'd356	:	dt	<=	92	;
						10'd357	:	dt	<=	92	;
						10'd358	:	dt	<=	144	;
						10'd359	:	dt	<=	241	;
						10'd360	:	dt	<=	231	;
						10'd361	:	dt	<=	233	;
						10'd362	:	dt	<=	233	;
						10'd363	:	dt	<=	234	;
						10'd364	:	dt	<=	206	;
						10'd365	:	dt	<=	209	;
						10'd366	:	dt	<=	211	;
						10'd367	:	dt	<=	214	;
						10'd368	:	dt	<=	228	;
						10'd369	:	dt	<=	218	;
						10'd370	:	dt	<=	196	;
						10'd371	:	dt	<=	186	;
						10'd372	:	dt	<=	171	;
						10'd373	:	dt	<=	116	;
						10'd374	:	dt	<=	162	;
						10'd375	:	dt	<=	161	;
						10'd376	:	dt	<=	123	;
						10'd377	:	dt	<=	50	;
						10'd378	:	dt	<=	205	;
						10'd379	:	dt	<=	255	;
						10'd380	:	dt	<=	203	;
						10'd381	:	dt	<=	153	;
						10'd382	:	dt	<=	111	;
						10'd383	:	dt	<=	97	;
						10'd384	:	dt	<=	98	;
						10'd385	:	dt	<=	96	;
						10'd386	:	dt	<=	162	;
						10'd387	:	dt	<=	244	;
						10'd388	:	dt	<=	228	;
						10'd389	:	dt	<=	233	;
						10'd390	:	dt	<=	233	;
						10'd391	:	dt	<=	235	;
						10'd392	:	dt	<=	208	;
						10'd393	:	dt	<=	209	;
						10'd394	:	dt	<=	208	;
						10'd395	:	dt	<=	225	;
						10'd396	:	dt	<=	241	;
						10'd397	:	dt	<=	203	;
						10'd398	:	dt	<=	187	;
						10'd399	:	dt	<=	156	;
						10'd400	:	dt	<=	136	;
						10'd401	:	dt	<=	102	;
						10'd402	:	dt	<=	131	;
						10'd403	:	dt	<=	147	;
						10'd404	:	dt	<=	89	;
						10'd405	:	dt	<=	105	;
						10'd406	:	dt	<=	255	;
						10'd407	:	dt	<=	239	;
						10'd408	:	dt	<=	198	;
						10'd409	:	dt	<=	156	;
						10'd410	:	dt	<=	115	;
						10'd411	:	dt	<=	90	;
						10'd412	:	dt	<=	98	;
						10'd413	:	dt	<=	96	;
						10'd414	:	dt	<=	178	;
						10'd415	:	dt	<=	245	;
						10'd416	:	dt	<=	232	;
						10'd417	:	dt	<=	235	;
						10'd418	:	dt	<=	235	;
						10'd419	:	dt	<=	235	;
						10'd420	:	dt	<=	208	;
						10'd421	:	dt	<=	211	;
						10'd422	:	dt	<=	209	;
						10'd423	:	dt	<=	227	;
						10'd424	:	dt	<=	251	;
						10'd425	:	dt	<=	217	;
						10'd426	:	dt	<=	192	;
						10'd427	:	dt	<=	164	;
						10'd428	:	dt	<=	159	;
						10'd429	:	dt	<=	105	;
						10'd430	:	dt	<=	131	;
						10'd431	:	dt	<=	148	;
						10'd432	:	dt	<=	167	;
						10'd433	:	dt	<=	239	;
						10'd434	:	dt	<=	255	;
						10'd435	:	dt	<=	229	;
						10'd436	:	dt	<=	192	;
						10'd437	:	dt	<=	156	;
						10'd438	:	dt	<=	118	;
						10'd439	:	dt	<=	101	;
						10'd440	:	dt	<=	104	;
						10'd441	:	dt	<=	107	;
						10'd442	:	dt	<=	218	;
						10'd443	:	dt	<=	238	;
						10'd444	:	dt	<=	234	;
						10'd445	:	dt	<=	236	;
						10'd446	:	dt	<=	236	;
						10'd447	:	dt	<=	236	;
						10'd448	:	dt	<=	209	;
						10'd449	:	dt	<=	213	;
						10'd450	:	dt	<=	206	;
						10'd451	:	dt	<=	240	;
						10'd452	:	dt	<=	247	;
						10'd453	:	dt	<=	214	;
						10'd454	:	dt	<=	192	;
						10'd455	:	dt	<=	169	;
						10'd456	:	dt	<=	160	;
						10'd457	:	dt	<=	139	;
						10'd458	:	dt	<=	145	;
						10'd459	:	dt	<=	205	;
						10'd460	:	dt	<=	255	;
						10'd461	:	dt	<=	240	;
						10'd462	:	dt	<=	224	;
						10'd463	:	dt	<=	218	;
						10'd464	:	dt	<=	186	;
						10'd465	:	dt	<=	146	;
						10'd466	:	dt	<=	114	;
						10'd467	:	dt	<=	105	;
						10'd468	:	dt	<=	92	;
						10'd469	:	dt	<=	133	;
						10'd470	:	dt	<=	244	;
						10'd471	:	dt	<=	232	;
						10'd472	:	dt	<=	235	;
						10'd473	:	dt	<=	235	;
						10'd474	:	dt	<=	235	;
						10'd475	:	dt	<=	234	;
						10'd476	:	dt	<=	211	;
						10'd477	:	dt	<=	210	;
						10'd478	:	dt	<=	210	;
						10'd479	:	dt	<=	255	;
						10'd480	:	dt	<=	238	;
						10'd481	:	dt	<=	214	;
						10'd482	:	dt	<=	192	;
						10'd483	:	dt	<=	173	;
						10'd484	:	dt	<=	170	;
						10'd485	:	dt	<=	172	;
						10'd486	:	dt	<=	194	;
						10'd487	:	dt	<=	255	;
						10'd488	:	dt	<=	255	;
						10'd489	:	dt	<=	232	;
						10'd490	:	dt	<=	202	;
						10'd491	:	dt	<=	202	;
						10'd492	:	dt	<=	174	;
						10'd493	:	dt	<=	132	;
						10'd494	:	dt	<=	110	;
						10'd495	:	dt	<=	109	;
						10'd496	:	dt	<=	103	;
						10'd497	:	dt	<=	203	;
						10'd498	:	dt	<=	240	;
						10'd499	:	dt	<=	233	;
						10'd500	:	dt	<=	233	;
						10'd501	:	dt	<=	234	;
						10'd502	:	dt	<=	233	;
						10'd503	:	dt	<=	231	;
						10'd504	:	dt	<=	211	;
						10'd505	:	dt	<=	208	;
						10'd506	:	dt	<=	221	;
						10'd507	:	dt	<=	255	;
						10'd508	:	dt	<=	232	;
						10'd509	:	dt	<=	214	;
						10'd510	:	dt	<=	204	;
						10'd511	:	dt	<=	183	;
						10'd512	:	dt	<=	180	;
						10'd513	:	dt	<=	175	;
						10'd514	:	dt	<=	247	;
						10'd515	:	dt	<=	255	;
						10'd516	:	dt	<=	253	;
						10'd517	:	dt	<=	223	;
						10'd518	:	dt	<=	187	;
						10'd519	:	dt	<=	186	;
						10'd520	:	dt	<=	162	;
						10'd521	:	dt	<=	120	;
						10'd522	:	dt	<=	114	;
						10'd523	:	dt	<=	103	;
						10'd524	:	dt	<=	184	;
						10'd525	:	dt	<=	242	;
						10'd526	:	dt	<=	232	;
						10'd527	:	dt	<=	235	;
						10'd528	:	dt	<=	234	;
						10'd529	:	dt	<=	234	;
						10'd530	:	dt	<=	233	;
						10'd531	:	dt	<=	232	;
						10'd532	:	dt	<=	212	;
						10'd533	:	dt	<=	207	;
						10'd534	:	dt	<=	231	;
						10'd535	:	dt	<=	255	;
						10'd536	:	dt	<=	231	;
						10'd537	:	dt	<=	223	;
						10'd538	:	dt	<=	214	;
						10'd539	:	dt	<=	184	;
						10'd540	:	dt	<=	186	;
						10'd541	:	dt	<=	222	;
						10'd542	:	dt	<=	255	;
						10'd543	:	dt	<=	255	;
						10'd544	:	dt	<=	240	;
						10'd545	:	dt	<=	214	;
						10'd546	:	dt	<=	178	;
						10'd547	:	dt	<=	171	;
						10'd548	:	dt	<=	151	;
						10'd549	:	dt	<=	117	;
						10'd550	:	dt	<=	102	;
						10'd551	:	dt	<=	153	;
						10'd552	:	dt	<=	244	;
						10'd553	:	dt	<=	233	;
						10'd554	:	dt	<=	235	;
						10'd555	:	dt	<=	235	;
						10'd556	:	dt	<=	236	;
						10'd557	:	dt	<=	235	;
						10'd558	:	dt	<=	234	;
						10'd559	:	dt	<=	234	;
						10'd560	:	dt	<=	212	;
						10'd561	:	dt	<=	208	;
						10'd562	:	dt	<=	233	;
						10'd563	:	dt	<=	255	;
						10'd564	:	dt	<=	235	;
						10'd565	:	dt	<=	228	;
						10'd566	:	dt	<=	218	;
						10'd567	:	dt	<=	186	;
						10'd568	:	dt	<=	209	;
						10'd569	:	dt	<=	254	;
						10'd570	:	dt	<=	255	;
						10'd571	:	dt	<=	250	;
						10'd572	:	dt	<=	232	;
						10'd573	:	dt	<=	198	;
						10'd574	:	dt	<=	170	;
						10'd575	:	dt	<=	159	;
						10'd576	:	dt	<=	138	;
						10'd577	:	dt	<=	108	;
						10'd578	:	dt	<=	115	;
						10'd579	:	dt	<=	228	;
						10'd580	:	dt	<=	237	;
						10'd581	:	dt	<=	235	;
						10'd582	:	dt	<=	235	;
						10'd583	:	dt	<=	235	;
						10'd584	:	dt	<=	236	;
						10'd585	:	dt	<=	236	;
						10'd586	:	dt	<=	235	;
						10'd587	:	dt	<=	235	;
						10'd588	:	dt	<=	212	;
						10'd589	:	dt	<=	210	;
						10'd590	:	dt	<=	227	;
						10'd591	:	dt	<=	255	;
						10'd592	:	dt	<=	239	;
						10'd593	:	dt	<=	232	;
						10'd594	:	dt	<=	218	;
						10'd595	:	dt	<=	196	;
						10'd596	:	dt	<=	223	;
						10'd597	:	dt	<=	253	;
						10'd598	:	dt	<=	244	;
						10'd599	:	dt	<=	229	;
						10'd600	:	dt	<=	226	;
						10'd601	:	dt	<=	185	;
						10'd602	:	dt	<=	162	;
						10'd603	:	dt	<=	148	;
						10'd604	:	dt	<=	127	;
						10'd605	:	dt	<=	97	;
						10'd606	:	dt	<=	181	;
						10'd607	:	dt	<=	244	;
						10'd608	:	dt	<=	234	;
						10'd609	:	dt	<=	236	;
						10'd610	:	dt	<=	235	;
						10'd611	:	dt	<=	236	;
						10'd612	:	dt	<=	236	;
						10'd613	:	dt	<=	236	;
						10'd614	:	dt	<=	236	;
						10'd615	:	dt	<=	235	;
						10'd616	:	dt	<=	213	;
						10'd617	:	dt	<=	210	;
						10'd618	:	dt	<=	224	;
						10'd619	:	dt	<=	255	;
						10'd620	:	dt	<=	241	;
						10'd621	:	dt	<=	230	;
						10'd622	:	dt	<=	215	;
						10'd623	:	dt	<=	211	;
						10'd624	:	dt	<=	222	;
						10'd625	:	dt	<=	248	;
						10'd626	:	dt	<=	229	;
						10'd627	:	dt	<=	221	;
						10'd628	:	dt	<=	201	;
						10'd629	:	dt	<=	181	;
						10'd630	:	dt	<=	149	;
						10'd631	:	dt	<=	138	;
						10'd632	:	dt	<=	114	;
						10'd633	:	dt	<=	121	;
						10'd634	:	dt	<=	236	;
						10'd635	:	dt	<=	234	;
						10'd636	:	dt	<=	236	;
						10'd637	:	dt	<=	236	;
						10'd638	:	dt	<=	236	;
						10'd639	:	dt	<=	237	;
						10'd640	:	dt	<=	238	;
						10'd641	:	dt	<=	236	;
						10'd642	:	dt	<=	234	;
						10'd643	:	dt	<=	236	;
						10'd644	:	dt	<=	214	;
						10'd645	:	dt	<=	208	;
						10'd646	:	dt	<=	229	;
						10'd647	:	dt	<=	253	;
						10'd648	:	dt	<=	233	;
						10'd649	:	dt	<=	222	;
						10'd650	:	dt	<=	211	;
						10'd651	:	dt	<=	216	;
						10'd652	:	dt	<=	221	;
						10'd653	:	dt	<=	237	;
						10'd654	:	dt	<=	215	;
						10'd655	:	dt	<=	217	;
						10'd656	:	dt	<=	184	;
						10'd657	:	dt	<=	174	;
						10'd658	:	dt	<=	139	;
						10'd659	:	dt	<=	129	;
						10'd660	:	dt	<=	97	;
						10'd661	:	dt	<=	171	;
						10'd662	:	dt	<=	248	;
						10'd663	:	dt	<=	234	;
						10'd664	:	dt	<=	236	;
						10'd665	:	dt	<=	237	;
						10'd666	:	dt	<=	237	;
						10'd667	:	dt	<=	238	;
						10'd668	:	dt	<=	238	;
						10'd669	:	dt	<=	237	;
						10'd670	:	dt	<=	235	;
						10'd671	:	dt	<=	234	;
						10'd672	:	dt	<=	213	;
						10'd673	:	dt	<=	208	;
						10'd674	:	dt	<=	236	;
						10'd675	:	dt	<=	236	;
						10'd676	:	dt	<=	218	;
						10'd677	:	dt	<=	215	;
						10'd678	:	dt	<=	208	;
						10'd679	:	dt	<=	215	;
						10'd680	:	dt	<=	225	;
						10'd681	:	dt	<=	224	;
						10'd682	:	dt	<=	202	;
						10'd683	:	dt	<=	215	;
						10'd684	:	dt	<=	196	;
						10'd685	:	dt	<=	156	;
						10'd686	:	dt	<=	134	;
						10'd687	:	dt	<=	121	;
						10'd688	:	dt	<=	101	;
						10'd689	:	dt	<=	216	;
						10'd690	:	dt	<=	239	;
						10'd691	:	dt	<=	235	;
						10'd692	:	dt	<=	236	;
						10'd693	:	dt	<=	236	;
						10'd694	:	dt	<=	237	;
						10'd695	:	dt	<=	238	;
						10'd696	:	dt	<=	238	;
						10'd697	:	dt	<=	238	;
						10'd698	:	dt	<=	236	;
						10'd699	:	dt	<=	235	;
						10'd700	:	dt	<=	213	;
						10'd701	:	dt	<=	209	;
						10'd702	:	dt	<=	238	;
						10'd703	:	dt	<=	216	;
						10'd704	:	dt	<=	207	;
						10'd705	:	dt	<=	212	;
						10'd706	:	dt	<=	209	;
						10'd707	:	dt	<=	212	;
						10'd708	:	dt	<=	225	;
						10'd709	:	dt	<=	216	;
						10'd710	:	dt	<=	202	;
						10'd711	:	dt	<=	215	;
						10'd712	:	dt	<=	195	;
						10'd713	:	dt	<=	149	;
						10'd714	:	dt	<=	128	;
						10'd715	:	dt	<=	103	;
						10'd716	:	dt	<=	147	;
						10'd717	:	dt	<=	246	;
						10'd718	:	dt	<=	231	;
						10'd719	:	dt	<=	236	;
						10'd720	:	dt	<=	237	;
						10'd721	:	dt	<=	236	;
						10'd722	:	dt	<=	236	;
						10'd723	:	dt	<=	237	;
						10'd724	:	dt	<=	238	;
						10'd725	:	dt	<=	236	;
						10'd726	:	dt	<=	236	;
						10'd727	:	dt	<=	236	;
						10'd728	:	dt	<=	212	;
						10'd729	:	dt	<=	209	;
						10'd730	:	dt	<=	248	;
						10'd731	:	dt	<=	230	;
						10'd732	:	dt	<=	219	;
						10'd733	:	dt	<=	220	;
						10'd734	:	dt	<=	223	;
						10'd735	:	dt	<=	221	;
						10'd736	:	dt	<=	230	;
						10'd737	:	dt	<=	208	;
						10'd738	:	dt	<=	198	;
						10'd739	:	dt	<=	203	;
						10'd740	:	dt	<=	177	;
						10'd741	:	dt	<=	142	;
						10'd742	:	dt	<=	117	;
						10'd743	:	dt	<=	113	;
						10'd744	:	dt	<=	222	;
						10'd745	:	dt	<=	238	;
						10'd746	:	dt	<=	236	;
						10'd747	:	dt	<=	238	;
						10'd748	:	dt	<=	237	;
						10'd749	:	dt	<=	237	;
						10'd750	:	dt	<=	238	;
						10'd751	:	dt	<=	238	;
						10'd752	:	dt	<=	239	;
						10'd753	:	dt	<=	237	;
						10'd754	:	dt	<=	236	;
						10'd755	:	dt	<=	237	;
						10'd756	:	dt	<=	210	;
						10'd757	:	dt	<=	213	;
						10'd758	:	dt	<=	255	;
						10'd759	:	dt	<=	241	;
						10'd760	:	dt	<=	221	;
						10'd761	:	dt	<=	225	;
						10'd762	:	dt	<=	232	;
						10'd763	:	dt	<=	226	;
						10'd764	:	dt	<=	234	;
						10'd765	:	dt	<=	190	;
						10'd766	:	dt	<=	188	;
						10'd767	:	dt	<=	188	;
						10'd768	:	dt	<=	158	;
						10'd769	:	dt	<=	133	;
						10'd770	:	dt	<=	103	;
						10'd771	:	dt	<=	188	;
						10'd772	:	dt	<=	246	;
						10'd773	:	dt	<=	235	;
						10'd774	:	dt	<=	237	;
						10'd775	:	dt	<=	237	;
						10'd776	:	dt	<=	238	;
						10'd777	:	dt	<=	239	;
						10'd778	:	dt	<=	239	;
						10'd779	:	dt	<=	239	;
						10'd780	:	dt	<=	239	;
						10'd781	:	dt	<=	238	;
						10'd782	:	dt	<=	237	;
						10'd783	:	dt	<=	237	;
					endcase
				end
				5'd19	:	begin
					case (cnt)	
						10'd0	:	dt	<=	143	;
						10'd1	:	dt	<=	145	;
						10'd2	:	dt	<=	148	;
						10'd3	:	dt	<=	150	;
						10'd4	:	dt	<=	151	;
						10'd5	:	dt	<=	154	;
						10'd6	:	dt	<=	155	;
						10'd7	:	dt	<=	156	;
						10'd8	:	dt	<=	157	;
						10'd9	:	dt	<=	158	;
						10'd10	:	dt	<=	158	;
						10'd11	:	dt	<=	158	;
						10'd12	:	dt	<=	159	;
						10'd13	:	dt	<=	160	;
						10'd14	:	dt	<=	161	;
						10'd15	:	dt	<=	161	;
						10'd16	:	dt	<=	161	;
						10'd17	:	dt	<=	162	;
						10'd18	:	dt	<=	162	;
						10'd19	:	dt	<=	161	;
						10'd20	:	dt	<=	162	;
						10'd21	:	dt	<=	161	;
						10'd22	:	dt	<=	162	;
						10'd23	:	dt	<=	162	;
						10'd24	:	dt	<=	161	;
						10'd25	:	dt	<=	160	;
						10'd26	:	dt	<=	161	;
						10'd27	:	dt	<=	159	;
						10'd28	:	dt	<=	145	;
						10'd29	:	dt	<=	147	;
						10'd30	:	dt	<=	151	;
						10'd31	:	dt	<=	154	;
						10'd32	:	dt	<=	155	;
						10'd33	:	dt	<=	157	;
						10'd34	:	dt	<=	159	;
						10'd35	:	dt	<=	160	;
						10'd36	:	dt	<=	160	;
						10'd37	:	dt	<=	161	;
						10'd38	:	dt	<=	160	;
						10'd39	:	dt	<=	161	;
						10'd40	:	dt	<=	162	;
						10'd41	:	dt	<=	164	;
						10'd42	:	dt	<=	165	;
						10'd43	:	dt	<=	165	;
						10'd44	:	dt	<=	164	;
						10'd45	:	dt	<=	164	;
						10'd46	:	dt	<=	164	;
						10'd47	:	dt	<=	165	;
						10'd48	:	dt	<=	165	;
						10'd49	:	dt	<=	164	;
						10'd50	:	dt	<=	165	;
						10'd51	:	dt	<=	165	;
						10'd52	:	dt	<=	164	;
						10'd53	:	dt	<=	164	;
						10'd54	:	dt	<=	164	;
						10'd55	:	dt	<=	162	;
						10'd56	:	dt	<=	149	;
						10'd57	:	dt	<=	151	;
						10'd58	:	dt	<=	155	;
						10'd59	:	dt	<=	158	;
						10'd60	:	dt	<=	160	;
						10'd61	:	dt	<=	161	;
						10'd62	:	dt	<=	162	;
						10'd63	:	dt	<=	164	;
						10'd64	:	dt	<=	164	;
						10'd65	:	dt	<=	165	;
						10'd66	:	dt	<=	165	;
						10'd67	:	dt	<=	165	;
						10'd68	:	dt	<=	165	;
						10'd69	:	dt	<=	165	;
						10'd70	:	dt	<=	167	;
						10'd71	:	dt	<=	167	;
						10'd72	:	dt	<=	167	;
						10'd73	:	dt	<=	168	;
						10'd74	:	dt	<=	168	;
						10'd75	:	dt	<=	168	;
						10'd76	:	dt	<=	168	;
						10'd77	:	dt	<=	167	;
						10'd78	:	dt	<=	167	;
						10'd79	:	dt	<=	167	;
						10'd80	:	dt	<=	166	;
						10'd81	:	dt	<=	167	;
						10'd82	:	dt	<=	166	;
						10'd83	:	dt	<=	165	;
						10'd84	:	dt	<=	153	;
						10'd85	:	dt	<=	155	;
						10'd86	:	dt	<=	159	;
						10'd87	:	dt	<=	162	;
						10'd88	:	dt	<=	163	;
						10'd89	:	dt	<=	164	;
						10'd90	:	dt	<=	165	;
						10'd91	:	dt	<=	166	;
						10'd92	:	dt	<=	167	;
						10'd93	:	dt	<=	168	;
						10'd94	:	dt	<=	168	;
						10'd95	:	dt	<=	171	;
						10'd96	:	dt	<=	164	;
						10'd97	:	dt	<=	134	;
						10'd98	:	dt	<=	143	;
						10'd99	:	dt	<=	171	;
						10'd100	:	dt	<=	170	;
						10'd101	:	dt	<=	171	;
						10'd102	:	dt	<=	172	;
						10'd103	:	dt	<=	172	;
						10'd104	:	dt	<=	172	;
						10'd105	:	dt	<=	171	;
						10'd106	:	dt	<=	171	;
						10'd107	:	dt	<=	171	;
						10'd108	:	dt	<=	170	;
						10'd109	:	dt	<=	170	;
						10'd110	:	dt	<=	169	;
						10'd111	:	dt	<=	167	;
						10'd112	:	dt	<=	156	;
						10'd113	:	dt	<=	158	;
						10'd114	:	dt	<=	162	;
						10'd115	:	dt	<=	164	;
						10'd116	:	dt	<=	166	;
						10'd117	:	dt	<=	167	;
						10'd118	:	dt	<=	167	;
						10'd119	:	dt	<=	169	;
						10'd120	:	dt	<=	170	;
						10'd121	:	dt	<=	171	;
						10'd122	:	dt	<=	171	;
						10'd123	:	dt	<=	180	;
						10'd124	:	dt	<=	169	;
						10'd125	:	dt	<=	132	;
						10'd126	:	dt	<=	100	;
						10'd127	:	dt	<=	172	;
						10'd128	:	dt	<=	174	;
						10'd129	:	dt	<=	175	;
						10'd130	:	dt	<=	174	;
						10'd131	:	dt	<=	174	;
						10'd132	:	dt	<=	174	;
						10'd133	:	dt	<=	173	;
						10'd134	:	dt	<=	174	;
						10'd135	:	dt	<=	175	;
						10'd136	:	dt	<=	174	;
						10'd137	:	dt	<=	174	;
						10'd138	:	dt	<=	173	;
						10'd139	:	dt	<=	172	;
						10'd140	:	dt	<=	158	;
						10'd141	:	dt	<=	161	;
						10'd142	:	dt	<=	164	;
						10'd143	:	dt	<=	167	;
						10'd144	:	dt	<=	169	;
						10'd145	:	dt	<=	171	;
						10'd146	:	dt	<=	171	;
						10'd147	:	dt	<=	172	;
						10'd148	:	dt	<=	173	;
						10'd149	:	dt	<=	173	;
						10'd150	:	dt	<=	175	;
						10'd151	:	dt	<=	185	;
						10'd152	:	dt	<=	174	;
						10'd153	:	dt	<=	136	;
						10'd154	:	dt	<=	86	;
						10'd155	:	dt	<=	163	;
						10'd156	:	dt	<=	178	;
						10'd157	:	dt	<=	178	;
						10'd158	:	dt	<=	179	;
						10'd159	:	dt	<=	178	;
						10'd160	:	dt	<=	177	;
						10'd161	:	dt	<=	177	;
						10'd162	:	dt	<=	177	;
						10'd163	:	dt	<=	177	;
						10'd164	:	dt	<=	177	;
						10'd165	:	dt	<=	177	;
						10'd166	:	dt	<=	176	;
						10'd167	:	dt	<=	175	;
						10'd168	:	dt	<=	161	;
						10'd169	:	dt	<=	165	;
						10'd170	:	dt	<=	167	;
						10'd171	:	dt	<=	170	;
						10'd172	:	dt	<=	172	;
						10'd173	:	dt	<=	174	;
						10'd174	:	dt	<=	174	;
						10'd175	:	dt	<=	176	;
						10'd176	:	dt	<=	177	;
						10'd177	:	dt	<=	178	;
						10'd178	:	dt	<=	179	;
						10'd179	:	dt	<=	185	;
						10'd180	:	dt	<=	175	;
						10'd181	:	dt	<=	137	;
						10'd182	:	dt	<=	91	;
						10'd183	:	dt	<=	146	;
						10'd184	:	dt	<=	157	;
						10'd185	:	dt	<=	161	;
						10'd186	:	dt	<=	175	;
						10'd187	:	dt	<=	177	;
						10'd188	:	dt	<=	177	;
						10'd189	:	dt	<=	180	;
						10'd190	:	dt	<=	180	;
						10'd191	:	dt	<=	180	;
						10'd192	:	dt	<=	180	;
						10'd193	:	dt	<=	180	;
						10'd194	:	dt	<=	179	;
						10'd195	:	dt	<=	178	;
						10'd196	:	dt	<=	165	;
						10'd197	:	dt	<=	168	;
						10'd198	:	dt	<=	170	;
						10'd199	:	dt	<=	172	;
						10'd200	:	dt	<=	174	;
						10'd201	:	dt	<=	175	;
						10'd202	:	dt	<=	177	;
						10'd203	:	dt	<=	178	;
						10'd204	:	dt	<=	181	;
						10'd205	:	dt	<=	182	;
						10'd206	:	dt	<=	182	;
						10'd207	:	dt	<=	183	;
						10'd208	:	dt	<=	169	;
						10'd209	:	dt	<=	155	;
						10'd210	:	dt	<=	158	;
						10'd211	:	dt	<=	165	;
						10'd212	:	dt	<=	148	;
						10'd213	:	dt	<=	121	;
						10'd214	:	dt	<=	140	;
						10'd215	:	dt	<=	143	;
						10'd216	:	dt	<=	140	;
						10'd217	:	dt	<=	148	;
						10'd218	:	dt	<=	153	;
						10'd219	:	dt	<=	173	;
						10'd220	:	dt	<=	173	;
						10'd221	:	dt	<=	179	;
						10'd222	:	dt	<=	181	;
						10'd223	:	dt	<=	179	;
						10'd224	:	dt	<=	167	;
						10'd225	:	dt	<=	170	;
						10'd226	:	dt	<=	173	;
						10'd227	:	dt	<=	175	;
						10'd228	:	dt	<=	177	;
						10'd229	:	dt	<=	179	;
						10'd230	:	dt	<=	180	;
						10'd231	:	dt	<=	181	;
						10'd232	:	dt	<=	178	;
						10'd233	:	dt	<=	175	;
						10'd234	:	dt	<=	175	;
						10'd235	:	dt	<=	174	;
						10'd236	:	dt	<=	174	;
						10'd237	:	dt	<=	173	;
						10'd238	:	dt	<=	167	;
						10'd239	:	dt	<=	157	;
						10'd240	:	dt	<=	140	;
						10'd241	:	dt	<=	113	;
						10'd242	:	dt	<=	125	;
						10'd243	:	dt	<=	143	;
						10'd244	:	dt	<=	143	;
						10'd245	:	dt	<=	141	;
						10'd246	:	dt	<=	131	;
						10'd247	:	dt	<=	149	;
						10'd248	:	dt	<=	141	;
						10'd249	:	dt	<=	167	;
						10'd250	:	dt	<=	184	;
						10'd251	:	dt	<=	183	;
						10'd252	:	dt	<=	170	;
						10'd253	:	dt	<=	173	;
						10'd254	:	dt	<=	175	;
						10'd255	:	dt	<=	178	;
						10'd256	:	dt	<=	180	;
						10'd257	:	dt	<=	181	;
						10'd258	:	dt	<=	182	;
						10'd259	:	dt	<=	177	;
						10'd260	:	dt	<=	154	;
						10'd261	:	dt	<=	153	;
						10'd262	:	dt	<=	158	;
						10'd263	:	dt	<=	160	;
						10'd264	:	dt	<=	160	;
						10'd265	:	dt	<=	157	;
						10'd266	:	dt	<=	153	;
						10'd267	:	dt	<=	155	;
						10'd268	:	dt	<=	145	;
						10'd269	:	dt	<=	112	;
						10'd270	:	dt	<=	97	;
						10'd271	:	dt	<=	115	;
						10'd272	:	dt	<=	122	;
						10'd273	:	dt	<=	118	;
						10'd274	:	dt	<=	114	;
						10'd275	:	dt	<=	117	;
						10'd276	:	dt	<=	141	;
						10'd277	:	dt	<=	181	;
						10'd278	:	dt	<=	186	;
						10'd279	:	dt	<=	185	;
						10'd280	:	dt	<=	172	;
						10'd281	:	dt	<=	175	;
						10'd282	:	dt	<=	177	;
						10'd283	:	dt	<=	180	;
						10'd284	:	dt	<=	182	;
						10'd285	:	dt	<=	184	;
						10'd286	:	dt	<=	186	;
						10'd287	:	dt	<=	167	;
						10'd288	:	dt	<=	146	;
						10'd289	:	dt	<=	142	;
						10'd290	:	dt	<=	141	;
						10'd291	:	dt	<=	147	;
						10'd292	:	dt	<=	151	;
						10'd293	:	dt	<=	155	;
						10'd294	:	dt	<=	153	;
						10'd295	:	dt	<=	153	;
						10'd296	:	dt	<=	143	;
						10'd297	:	dt	<=	104	;
						10'd298	:	dt	<=	155	;
						10'd299	:	dt	<=	176	;
						10'd300	:	dt	<=	176	;
						10'd301	:	dt	<=	169	;
						10'd302	:	dt	<=	172	;
						10'd303	:	dt	<=	177	;
						10'd304	:	dt	<=	187	;
						10'd305	:	dt	<=	189	;
						10'd306	:	dt	<=	188	;
						10'd307	:	dt	<=	187	;
						10'd308	:	dt	<=	173	;
						10'd309	:	dt	<=	177	;
						10'd310	:	dt	<=	179	;
						10'd311	:	dt	<=	182	;
						10'd312	:	dt	<=	184	;
						10'd313	:	dt	<=	185	;
						10'd314	:	dt	<=	190	;
						10'd315	:	dt	<=	165	;
						10'd316	:	dt	<=	160	;
						10'd317	:	dt	<=	144	;
						10'd318	:	dt	<=	132	;
						10'd319	:	dt	<=	133	;
						10'd320	:	dt	<=	139	;
						10'd321	:	dt	<=	143	;
						10'd322	:	dt	<=	140	;
						10'd323	:	dt	<=	136	;
						10'd324	:	dt	<=	131	;
						10'd325	:	dt	<=	108	;
						10'd326	:	dt	<=	163	;
						10'd327	:	dt	<=	194	;
						10'd328	:	dt	<=	193	;
						10'd329	:	dt	<=	193	;
						10'd330	:	dt	<=	194	;
						10'd331	:	dt	<=	193	;
						10'd332	:	dt	<=	193	;
						10'd333	:	dt	<=	193	;
						10'd334	:	dt	<=	190	;
						10'd335	:	dt	<=	189	;
						10'd336	:	dt	<=	176	;
						10'd337	:	dt	<=	179	;
						10'd338	:	dt	<=	181	;
						10'd339	:	dt	<=	184	;
						10'd340	:	dt	<=	187	;
						10'd341	:	dt	<=	187	;
						10'd342	:	dt	<=	188	;
						10'd343	:	dt	<=	186	;
						10'd344	:	dt	<=	181	;
						10'd345	:	dt	<=	150	;
						10'd346	:	dt	<=	126	;
						10'd347	:	dt	<=	128	;
						10'd348	:	dt	<=	133	;
						10'd349	:	dt	<=	142	;
						10'd350	:	dt	<=	148	;
						10'd351	:	dt	<=	142	;
						10'd352	:	dt	<=	131	;
						10'd353	:	dt	<=	114	;
						10'd354	:	dt	<=	129	;
						10'd355	:	dt	<=	197	;
						10'd356	:	dt	<=	195	;
						10'd357	:	dt	<=	195	;
						10'd358	:	dt	<=	195	;
						10'd359	:	dt	<=	196	;
						10'd360	:	dt	<=	195	;
						10'd361	:	dt	<=	194	;
						10'd362	:	dt	<=	193	;
						10'd363	:	dt	<=	192	;
						10'd364	:	dt	<=	178	;
						10'd365	:	dt	<=	181	;
						10'd366	:	dt	<=	183	;
						10'd367	:	dt	<=	186	;
						10'd368	:	dt	<=	188	;
						10'd369	:	dt	<=	189	;
						10'd370	:	dt	<=	186	;
						10'd371	:	dt	<=	190	;
						10'd372	:	dt	<=	190	;
						10'd373	:	dt	<=	166	;
						10'd374	:	dt	<=	140	;
						10'd375	:	dt	<=	117	;
						10'd376	:	dt	<=	118	;
						10'd377	:	dt	<=	127	;
						10'd378	:	dt	<=	132	;
						10'd379	:	dt	<=	123	;
						10'd380	:	dt	<=	114	;
						10'd381	:	dt	<=	100	;
						10'd382	:	dt	<=	133	;
						10'd383	:	dt	<=	197	;
						10'd384	:	dt	<=	196	;
						10'd385	:	dt	<=	197	;
						10'd386	:	dt	<=	196	;
						10'd387	:	dt	<=	197	;
						10'd388	:	dt	<=	196	;
						10'd389	:	dt	<=	195	;
						10'd390	:	dt	<=	195	;
						10'd391	:	dt	<=	194	;
						10'd392	:	dt	<=	179	;
						10'd393	:	dt	<=	182	;
						10'd394	:	dt	<=	185	;
						10'd395	:	dt	<=	188	;
						10'd396	:	dt	<=	189	;
						10'd397	:	dt	<=	191	;
						10'd398	:	dt	<=	187	;
						10'd399	:	dt	<=	183	;
						10'd400	:	dt	<=	190	;
						10'd401	:	dt	<=	191	;
						10'd402	:	dt	<=	154	;
						10'd403	:	dt	<=	125	;
						10'd404	:	dt	<=	121	;
						10'd405	:	dt	<=	127	;
						10'd406	:	dt	<=	128	;
						10'd407	:	dt	<=	115	;
						10'd408	:	dt	<=	103	;
						10'd409	:	dt	<=	90	;
						10'd410	:	dt	<=	161	;
						10'd411	:	dt	<=	200	;
						10'd412	:	dt	<=	201	;
						10'd413	:	dt	<=	201	;
						10'd414	:	dt	<=	200	;
						10'd415	:	dt	<=	199	;
						10'd416	:	dt	<=	199	;
						10'd417	:	dt	<=	197	;
						10'd418	:	dt	<=	196	;
						10'd419	:	dt	<=	195	;
						10'd420	:	dt	<=	180	;
						10'd421	:	dt	<=	183	;
						10'd422	:	dt	<=	187	;
						10'd423	:	dt	<=	190	;
						10'd424	:	dt	<=	192	;
						10'd425	:	dt	<=	192	;
						10'd426	:	dt	<=	187	;
						10'd427	:	dt	<=	190	;
						10'd428	:	dt	<=	190	;
						10'd429	:	dt	<=	179	;
						10'd430	:	dt	<=	144	;
						10'd431	:	dt	<=	131	;
						10'd432	:	dt	<=	127	;
						10'd433	:	dt	<=	123	;
						10'd434	:	dt	<=	114	;
						10'd435	:	dt	<=	99	;
						10'd436	:	dt	<=	89	;
						10'd437	:	dt	<=	85	;
						10'd438	:	dt	<=	180	;
						10'd439	:	dt	<=	202	;
						10'd440	:	dt	<=	204	;
						10'd441	:	dt	<=	202	;
						10'd442	:	dt	<=	200	;
						10'd443	:	dt	<=	201	;
						10'd444	:	dt	<=	200	;
						10'd445	:	dt	<=	199	;
						10'd446	:	dt	<=	198	;
						10'd447	:	dt	<=	199	;
						10'd448	:	dt	<=	183	;
						10'd449	:	dt	<=	185	;
						10'd450	:	dt	<=	189	;
						10'd451	:	dt	<=	192	;
						10'd452	:	dt	<=	194	;
						10'd453	:	dt	<=	193	;
						10'd454	:	dt	<=	189	;
						10'd455	:	dt	<=	195	;
						10'd456	:	dt	<=	190	;
						10'd457	:	dt	<=	171	;
						10'd458	:	dt	<=	145	;
						10'd459	:	dt	<=	129	;
						10'd460	:	dt	<=	131	;
						10'd461	:	dt	<=	109	;
						10'd462	:	dt	<=	82	;
						10'd463	:	dt	<=	61	;
						10'd464	:	dt	<=	74	;
						10'd465	:	dt	<=	101	;
						10'd466	:	dt	<=	197	;
						10'd467	:	dt	<=	202	;
						10'd468	:	dt	<=	204	;
						10'd469	:	dt	<=	204	;
						10'd470	:	dt	<=	202	;
						10'd471	:	dt	<=	202	;
						10'd472	:	dt	<=	202	;
						10'd473	:	dt	<=	200	;
						10'd474	:	dt	<=	200	;
						10'd475	:	dt	<=	199	;
						10'd476	:	dt	<=	184	;
						10'd477	:	dt	<=	187	;
						10'd478	:	dt	<=	191	;
						10'd479	:	dt	<=	193	;
						10'd480	:	dt	<=	196	;
						10'd481	:	dt	<=	194	;
						10'd482	:	dt	<=	190	;
						10'd483	:	dt	<=	195	;
						10'd484	:	dt	<=	186	;
						10'd485	:	dt	<=	162	;
						10'd486	:	dt	<=	135	;
						10'd487	:	dt	<=	134	;
						10'd488	:	dt	<=	149	;
						10'd489	:	dt	<=	97	;
						10'd490	:	dt	<=	59	;
						10'd491	:	dt	<=	48	;
						10'd492	:	dt	<=	76	;
						10'd493	:	dt	<=	142	;
						10'd494	:	dt	<=	203	;
						10'd495	:	dt	<=	203	;
						10'd496	:	dt	<=	204	;
						10'd497	:	dt	<=	205	;
						10'd498	:	dt	<=	204	;
						10'd499	:	dt	<=	203	;
						10'd500	:	dt	<=	202	;
						10'd501	:	dt	<=	202	;
						10'd502	:	dt	<=	200	;
						10'd503	:	dt	<=	201	;
						10'd504	:	dt	<=	186	;
						10'd505	:	dt	<=	189	;
						10'd506	:	dt	<=	193	;
						10'd507	:	dt	<=	195	;
						10'd508	:	dt	<=	198	;
						10'd509	:	dt	<=	198	;
						10'd510	:	dt	<=	188	;
						10'd511	:	dt	<=	192	;
						10'd512	:	dt	<=	183	;
						10'd513	:	dt	<=	156	;
						10'd514	:	dt	<=	133	;
						10'd515	:	dt	<=	146	;
						10'd516	:	dt	<=	137	;
						10'd517	:	dt	<=	84	;
						10'd518	:	dt	<=	51	;
						10'd519	:	dt	<=	59	;
						10'd520	:	dt	<=	114	;
						10'd521	:	dt	<=	194	;
						10'd522	:	dt	<=	204	;
						10'd523	:	dt	<=	204	;
						10'd524	:	dt	<=	205	;
						10'd525	:	dt	<=	205	;
						10'd526	:	dt	<=	206	;
						10'd527	:	dt	<=	205	;
						10'd528	:	dt	<=	204	;
						10'd529	:	dt	<=	203	;
						10'd530	:	dt	<=	202	;
						10'd531	:	dt	<=	202	;
						10'd532	:	dt	<=	188	;
						10'd533	:	dt	<=	191	;
						10'd534	:	dt	<=	195	;
						10'd535	:	dt	<=	197	;
						10'd536	:	dt	<=	199	;
						10'd537	:	dt	<=	200	;
						10'd538	:	dt	<=	187	;
						10'd539	:	dt	<=	187	;
						10'd540	:	dt	<=	178	;
						10'd541	:	dt	<=	150	;
						10'd542	:	dt	<=	137	;
						10'd543	:	dt	<=	154	;
						10'd544	:	dt	<=	127	;
						10'd545	:	dt	<=	85	;
						10'd546	:	dt	<=	63	;
						10'd547	:	dt	<=	63	;
						10'd548	:	dt	<=	161	;
						10'd549	:	dt	<=	205	;
						10'd550	:	dt	<=	206	;
						10'd551	:	dt	<=	207	;
						10'd552	:	dt	<=	207	;
						10'd553	:	dt	<=	206	;
						10'd554	:	dt	<=	207	;
						10'd555	:	dt	<=	206	;
						10'd556	:	dt	<=	205	;
						10'd557	:	dt	<=	205	;
						10'd558	:	dt	<=	204	;
						10'd559	:	dt	<=	203	;
						10'd560	:	dt	<=	189	;
						10'd561	:	dt	<=	192	;
						10'd562	:	dt	<=	195	;
						10'd563	:	dt	<=	198	;
						10'd564	:	dt	<=	200	;
						10'd565	:	dt	<=	200	;
						10'd566	:	dt	<=	183	;
						10'd567	:	dt	<=	177	;
						10'd568	:	dt	<=	171	;
						10'd569	:	dt	<=	153	;
						10'd570	:	dt	<=	156	;
						10'd571	:	dt	<=	159	;
						10'd572	:	dt	<=	121	;
						10'd573	:	dt	<=	83	;
						10'd574	:	dt	<=	73	;
						10'd575	:	dt	<=	74	;
						10'd576	:	dt	<=	186	;
						10'd577	:	dt	<=	208	;
						10'd578	:	dt	<=	208	;
						10'd579	:	dt	<=	209	;
						10'd580	:	dt	<=	208	;
						10'd581	:	dt	<=	208	;
						10'd582	:	dt	<=	208	;
						10'd583	:	dt	<=	208	;
						10'd584	:	dt	<=	207	;
						10'd585	:	dt	<=	207	;
						10'd586	:	dt	<=	206	;
						10'd587	:	dt	<=	206	;
						10'd588	:	dt	<=	190	;
						10'd589	:	dt	<=	193	;
						10'd590	:	dt	<=	196	;
						10'd591	:	dt	<=	198	;
						10'd592	:	dt	<=	200	;
						10'd593	:	dt	<=	201	;
						10'd594	:	dt	<=	181	;
						10'd595	:	dt	<=	174	;
						10'd596	:	dt	<=	172	;
						10'd597	:	dt	<=	163	;
						10'd598	:	dt	<=	164	;
						10'd599	:	dt	<=	150	;
						10'd600	:	dt	<=	110	;
						10'd601	:	dt	<=	80	;
						10'd602	:	dt	<=	75	;
						10'd603	:	dt	<=	100	;
						10'd604	:	dt	<=	206	;
						10'd605	:	dt	<=	208	;
						10'd606	:	dt	<=	210	;
						10'd607	:	dt	<=	210	;
						10'd608	:	dt	<=	210	;
						10'd609	:	dt	<=	209	;
						10'd610	:	dt	<=	209	;
						10'd611	:	dt	<=	209	;
						10'd612	:	dt	<=	208	;
						10'd613	:	dt	<=	208	;
						10'd614	:	dt	<=	207	;
						10'd615	:	dt	<=	207	;
						10'd616	:	dt	<=	191	;
						10'd617	:	dt	<=	194	;
						10'd618	:	dt	<=	196	;
						10'd619	:	dt	<=	199	;
						10'd620	:	dt	<=	200	;
						10'd621	:	dt	<=	201	;
						10'd622	:	dt	<=	175	;
						10'd623	:	dt	<=	176	;
						10'd624	:	dt	<=	174	;
						10'd625	:	dt	<=	163	;
						10'd626	:	dt	<=	156	;
						10'd627	:	dt	<=	133	;
						10'd628	:	dt	<=	99	;
						10'd629	:	dt	<=	78	;
						10'd630	:	dt	<=	79	;
						10'd631	:	dt	<=	149	;
						10'd632	:	dt	<=	211	;
						10'd633	:	dt	<=	209	;
						10'd634	:	dt	<=	210	;
						10'd635	:	dt	<=	210	;
						10'd636	:	dt	<=	211	;
						10'd637	:	dt	<=	211	;
						10'd638	:	dt	<=	210	;
						10'd639	:	dt	<=	210	;
						10'd640	:	dt	<=	209	;
						10'd641	:	dt	<=	209	;
						10'd642	:	dt	<=	209	;
						10'd643	:	dt	<=	208	;
						10'd644	:	dt	<=	193	;
						10'd645	:	dt	<=	195	;
						10'd646	:	dt	<=	198	;
						10'd647	:	dt	<=	201	;
						10'd648	:	dt	<=	202	;
						10'd649	:	dt	<=	201	;
						10'd650	:	dt	<=	173	;
						10'd651	:	dt	<=	178	;
						10'd652	:	dt	<=	168	;
						10'd653	:	dt	<=	151	;
						10'd654	:	dt	<=	140	;
						10'd655	:	dt	<=	114	;
						10'd656	:	dt	<=	91	;
						10'd657	:	dt	<=	80	;
						10'd658	:	dt	<=	95	;
						10'd659	:	dt	<=	197	;
						10'd660	:	dt	<=	211	;
						10'd661	:	dt	<=	211	;
						10'd662	:	dt	<=	211	;
						10'd663	:	dt	<=	212	;
						10'd664	:	dt	<=	213	;
						10'd665	:	dt	<=	212	;
						10'd666	:	dt	<=	212	;
						10'd667	:	dt	<=	212	;
						10'd668	:	dt	<=	212	;
						10'd669	:	dt	<=	211	;
						10'd670	:	dt	<=	211	;
						10'd671	:	dt	<=	210	;
						10'd672	:	dt	<=	194	;
						10'd673	:	dt	<=	196	;
						10'd674	:	dt	<=	198	;
						10'd675	:	dt	<=	201	;
						10'd676	:	dt	<=	204	;
						10'd677	:	dt	<=	201	;
						10'd678	:	dt	<=	174	;
						10'd679	:	dt	<=	179	;
						10'd680	:	dt	<=	165	;
						10'd681	:	dt	<=	144	;
						10'd682	:	dt	<=	123	;
						10'd683	:	dt	<=	95	;
						10'd684	:	dt	<=	86	;
						10'd685	:	dt	<=	83	;
						10'd686	:	dt	<=	144	;
						10'd687	:	dt	<=	213	;
						10'd688	:	dt	<=	213	;
						10'd689	:	dt	<=	213	;
						10'd690	:	dt	<=	213	;
						10'd691	:	dt	<=	214	;
						10'd692	:	dt	<=	213	;
						10'd693	:	dt	<=	214	;
						10'd694	:	dt	<=	213	;
						10'd695	:	dt	<=	213	;
						10'd696	:	dt	<=	213	;
						10'd697	:	dt	<=	213	;
						10'd698	:	dt	<=	213	;
						10'd699	:	dt	<=	211	;
						10'd700	:	dt	<=	195	;
						10'd701	:	dt	<=	198	;
						10'd702	:	dt	<=	199	;
						10'd703	:	dt	<=	202	;
						10'd704	:	dt	<=	205	;
						10'd705	:	dt	<=	201	;
						10'd706	:	dt	<=	177	;
						10'd707	:	dt	<=	192	;
						10'd708	:	dt	<=	172	;
						10'd709	:	dt	<=	142	;
						10'd710	:	dt	<=	113	;
						10'd711	:	dt	<=	87	;
						10'd712	:	dt	<=	79	;
						10'd713	:	dt	<=	76	;
						10'd714	:	dt	<=	173	;
						10'd715	:	dt	<=	213	;
						10'd716	:	dt	<=	214	;
						10'd717	:	dt	<=	214	;
						10'd718	:	dt	<=	214	;
						10'd719	:	dt	<=	215	;
						10'd720	:	dt	<=	215	;
						10'd721	:	dt	<=	214	;
						10'd722	:	dt	<=	214	;
						10'd723	:	dt	<=	213	;
						10'd724	:	dt	<=	213	;
						10'd725	:	dt	<=	214	;
						10'd726	:	dt	<=	214	;
						10'd727	:	dt	<=	212	;
						10'd728	:	dt	<=	195	;
						10'd729	:	dt	<=	198	;
						10'd730	:	dt	<=	200	;
						10'd731	:	dt	<=	202	;
						10'd732	:	dt	<=	205	;
						10'd733	:	dt	<=	194	;
						10'd734	:	dt	<=	181	;
						10'd735	:	dt	<=	189	;
						10'd736	:	dt	<=	161	;
						10'd737	:	dt	<=	132	;
						10'd738	:	dt	<=	103	;
						10'd739	:	dt	<=	84	;
						10'd740	:	dt	<=	75	;
						10'd741	:	dt	<=	92	;
						10'd742	:	dt	<=	204	;
						10'd743	:	dt	<=	214	;
						10'd744	:	dt	<=	214	;
						10'd745	:	dt	<=	214	;
						10'd746	:	dt	<=	215	;
						10'd747	:	dt	<=	216	;
						10'd748	:	dt	<=	216	;
						10'd749	:	dt	<=	215	;
						10'd750	:	dt	<=	215	;
						10'd751	:	dt	<=	214	;
						10'd752	:	dt	<=	214	;
						10'd753	:	dt	<=	213	;
						10'd754	:	dt	<=	214	;
						10'd755	:	dt	<=	213	;
						10'd756	:	dt	<=	193	;
						10'd757	:	dt	<=	195	;
						10'd758	:	dt	<=	200	;
						10'd759	:	dt	<=	203	;
						10'd760	:	dt	<=	205	;
						10'd761	:	dt	<=	185	;
						10'd762	:	dt	<=	185	;
						10'd763	:	dt	<=	178	;
						10'd764	:	dt	<=	140	;
						10'd765	:	dt	<=	117	;
						10'd766	:	dt	<=	98	;
						10'd767	:	dt	<=	86	;
						10'd768	:	dt	<=	71	;
						10'd769	:	dt	<=	130	;
						10'd770	:	dt	<=	215	;
						10'd771	:	dt	<=	214	;
						10'd772	:	dt	<=	214	;
						10'd773	:	dt	<=	214	;
						10'd774	:	dt	<=	215	;
						10'd775	:	dt	<=	215	;
						10'd776	:	dt	<=	215	;
						10'd777	:	dt	<=	215	;
						10'd778	:	dt	<=	215	;
						10'd779	:	dt	<=	214	;
						10'd780	:	dt	<=	214	;
						10'd781	:	dt	<=	215	;
						10'd782	:	dt	<=	215	;
						10'd783	:	dt	<=	214	;				
					endcase
				end
				5'd20	:	begin
					case (cnt)
						10'd0	:	dt	<=	173	;
						10'd1	:	dt	<=	176	;
						10'd2	:	dt	<=	181	;
						10'd3	:	dt	<=	183	;
						10'd4	:	dt	<=	187	;
						10'd5	:	dt	<=	189	;
						10'd6	:	dt	<=	191	;
						10'd7	:	dt	<=	192	;
						10'd8	:	dt	<=	193	;
						10'd9	:	dt	<=	195	;
						10'd10	:	dt	<=	196	;
						10'd11	:	dt	<=	194	;
						10'd12	:	dt	<=	193	;
						10'd13	:	dt	<=	193	;
						10'd14	:	dt	<=	194	;
						10'd15	:	dt	<=	190	;
						10'd16	:	dt	<=	193	;
						10'd17	:	dt	<=	178	;
						10'd18	:	dt	<=	188	;
						10'd19	:	dt	<=	190	;
						10'd20	:	dt	<=	187	;
						10'd21	:	dt	<=	187	;
						10'd22	:	dt	<=	186	;
						10'd23	:	dt	<=	183	;
						10'd24	:	dt	<=	182	;
						10'd25	:	dt	<=	181	;
						10'd26	:	dt	<=	180	;
						10'd27	:	dt	<=	179	;
						10'd28	:	dt	<=	174	;
						10'd29	:	dt	<=	178	;
						10'd30	:	dt	<=	183	;
						10'd31	:	dt	<=	186	;
						10'd32	:	dt	<=	189	;
						10'd33	:	dt	<=	191	;
						10'd34	:	dt	<=	194	;
						10'd35	:	dt	<=	195	;
						10'd36	:	dt	<=	196	;
						10'd37	:	dt	<=	197	;
						10'd38	:	dt	<=	198	;
						10'd39	:	dt	<=	198	;
						10'd40	:	dt	<=	196	;
						10'd41	:	dt	<=	196	;
						10'd42	:	dt	<=	194	;
						10'd43	:	dt	<=	197	;
						10'd44	:	dt	<=	209	;
						10'd45	:	dt	<=	137	;
						10'd46	:	dt	<=	152	;
						10'd47	:	dt	<=	194	;
						10'd48	:	dt	<=	190	;
						10'd49	:	dt	<=	187	;
						10'd50	:	dt	<=	187	;
						10'd51	:	dt	<=	185	;
						10'd52	:	dt	<=	184	;
						10'd53	:	dt	<=	185	;
						10'd54	:	dt	<=	182	;
						10'd55	:	dt	<=	181	;
						10'd56	:	dt	<=	175	;
						10'd57	:	dt	<=	180	;
						10'd58	:	dt	<=	183	;
						10'd59	:	dt	<=	187	;
						10'd60	:	dt	<=	190	;
						10'd61	:	dt	<=	193	;
						10'd62	:	dt	<=	195	;
						10'd63	:	dt	<=	196	;
						10'd64	:	dt	<=	197	;
						10'd65	:	dt	<=	198	;
						10'd66	:	dt	<=	199	;
						10'd67	:	dt	<=	198	;
						10'd68	:	dt	<=	197	;
						10'd69	:	dt	<=	197	;
						10'd70	:	dt	<=	195	;
						10'd71	:	dt	<=	205	;
						10'd72	:	dt	<=	210	;
						10'd73	:	dt	<=	132	;
						10'd74	:	dt	<=	115	;
						10'd75	:	dt	<=	168	;
						10'd76	:	dt	<=	147	;
						10'd77	:	dt	<=	190	;
						10'd78	:	dt	<=	188	;
						10'd79	:	dt	<=	187	;
						10'd80	:	dt	<=	187	;
						10'd81	:	dt	<=	186	;
						10'd82	:	dt	<=	184	;
						10'd83	:	dt	<=	182	;
						10'd84	:	dt	<=	178	;
						10'd85	:	dt	<=	182	;
						10'd86	:	dt	<=	185	;
						10'd87	:	dt	<=	188	;
						10'd88	:	dt	<=	192	;
						10'd89	:	dt	<=	195	;
						10'd90	:	dt	<=	196	;
						10'd91	:	dt	<=	199	;
						10'd92	:	dt	<=	200	;
						10'd93	:	dt	<=	200	;
						10'd94	:	dt	<=	201	;
						10'd95	:	dt	<=	199	;
						10'd96	:	dt	<=	199	;
						10'd97	:	dt	<=	199	;
						10'd98	:	dt	<=	195	;
						10'd99	:	dt	<=	210	;
						10'd100	:	dt	<=	203	;
						10'd101	:	dt	<=	125	;
						10'd102	:	dt	<=	120	;
						10'd103	:	dt	<=	180	;
						10'd104	:	dt	<=	104	;
						10'd105	:	dt	<=	176	;
						10'd106	:	dt	<=	195	;
						10'd107	:	dt	<=	189	;
						10'd108	:	dt	<=	189	;
						10'd109	:	dt	<=	187	;
						10'd110	:	dt	<=	186	;
						10'd111	:	dt	<=	185	;
						10'd112	:	dt	<=	180	;
						10'd113	:	dt	<=	183	;
						10'd114	:	dt	<=	188	;
						10'd115	:	dt	<=	191	;
						10'd116	:	dt	<=	194	;
						10'd117	:	dt	<=	196	;
						10'd118	:	dt	<=	198	;
						10'd119	:	dt	<=	202	;
						10'd120	:	dt	<=	203	;
						10'd121	:	dt	<=	201	;
						10'd122	:	dt	<=	203	;
						10'd123	:	dt	<=	204	;
						10'd124	:	dt	<=	202	;
						10'd125	:	dt	<=	201	;
						10'd126	:	dt	<=	196	;
						10'd127	:	dt	<=	222	;
						10'd128	:	dt	<=	210	;
						10'd129	:	dt	<=	128	;
						10'd130	:	dt	<=	125	;
						10'd131	:	dt	<=	181	;
						10'd132	:	dt	<=	108	;
						10'd133	:	dt	<=	165	;
						10'd134	:	dt	<=	198	;
						10'd135	:	dt	<=	191	;
						10'd136	:	dt	<=	192	;
						10'd137	:	dt	<=	189	;
						10'd138	:	dt	<=	188	;
						10'd139	:	dt	<=	187	;
						10'd140	:	dt	<=	181	;
						10'd141	:	dt	<=	186	;
						10'd142	:	dt	<=	188	;
						10'd143	:	dt	<=	191	;
						10'd144	:	dt	<=	195	;
						10'd145	:	dt	<=	198	;
						10'd146	:	dt	<=	200	;
						10'd147	:	dt	<=	203	;
						10'd148	:	dt	<=	203	;
						10'd149	:	dt	<=	202	;
						10'd150	:	dt	<=	204	;
						10'd151	:	dt	<=	205	;
						10'd152	:	dt	<=	204	;
						10'd153	:	dt	<=	204	;
						10'd154	:	dt	<=	199	;
						10'd155	:	dt	<=	231	;
						10'd156	:	dt	<=	203	;
						10'd157	:	dt	<=	127	;
						10'd158	:	dt	<=	135	;
						10'd159	:	dt	<=	182	;
						10'd160	:	dt	<=	116	;
						10'd161	:	dt	<=	166	;
						10'd162	:	dt	<=	201	;
						10'd163	:	dt	<=	192	;
						10'd164	:	dt	<=	193	;
						10'd165	:	dt	<=	191	;
						10'd166	:	dt	<=	190	;
						10'd167	:	dt	<=	187	;
						10'd168	:	dt	<=	183	;
						10'd169	:	dt	<=	188	;
						10'd170	:	dt	<=	190	;
						10'd171	:	dt	<=	194	;
						10'd172	:	dt	<=	196	;
						10'd173	:	dt	<=	199	;
						10'd174	:	dt	<=	202	;
						10'd175	:	dt	<=	203	;
						10'd176	:	dt	<=	203	;
						10'd177	:	dt	<=	205	;
						10'd178	:	dt	<=	205	;
						10'd179	:	dt	<=	205	;
						10'd180	:	dt	<=	205	;
						10'd181	:	dt	<=	203	;
						10'd182	:	dt	<=	207	;
						10'd183	:	dt	<=	223	;
						10'd184	:	dt	<=	177	;
						10'd185	:	dt	<=	114	;
						10'd186	:	dt	<=	165	;
						10'd187	:	dt	<=	196	;
						10'd188	:	dt	<=	124	;
						10'd189	:	dt	<=	159	;
						10'd190	:	dt	<=	204	;
						10'd191	:	dt	<=	194	;
						10'd192	:	dt	<=	194	;
						10'd193	:	dt	<=	193	;
						10'd194	:	dt	<=	190	;
						10'd195	:	dt	<=	189	;
						10'd196	:	dt	<=	185	;
						10'd197	:	dt	<=	190	;
						10'd198	:	dt	<=	193	;
						10'd199	:	dt	<=	195	;
						10'd200	:	dt	<=	198	;
						10'd201	:	dt	<=	201	;
						10'd202	:	dt	<=	202	;
						10'd203	:	dt	<=	205	;
						10'd204	:	dt	<=	205	;
						10'd205	:	dt	<=	206	;
						10'd206	:	dt	<=	207	;
						10'd207	:	dt	<=	206	;
						10'd208	:	dt	<=	210	;
						10'd209	:	dt	<=	208	;
						10'd210	:	dt	<=	218	;
						10'd211	:	dt	<=	219	;
						10'd212	:	dt	<=	168	;
						10'd213	:	dt	<=	97	;
						10'd214	:	dt	<=	172	;
						10'd215	:	dt	<=	186	;
						10'd216	:	dt	<=	117	;
						10'd217	:	dt	<=	158	;
						10'd218	:	dt	<=	206	;
						10'd219	:	dt	<=	195	;
						10'd220	:	dt	<=	196	;
						10'd221	:	dt	<=	195	;
						10'd222	:	dt	<=	193	;
						10'd223	:	dt	<=	190	;
						10'd224	:	dt	<=	186	;
						10'd225	:	dt	<=	191	;
						10'd226	:	dt	<=	195	;
						10'd227	:	dt	<=	197	;
						10'd228	:	dt	<=	200	;
						10'd229	:	dt	<=	203	;
						10'd230	:	dt	<=	204	;
						10'd231	:	dt	<=	207	;
						10'd232	:	dt	<=	207	;
						10'd233	:	dt	<=	208	;
						10'd234	:	dt	<=	209	;
						10'd235	:	dt	<=	208	;
						10'd236	:	dt	<=	188	;
						10'd237	:	dt	<=	172	;
						10'd238	:	dt	<=	229	;
						10'd239	:	dt	<=	220	;
						10'd240	:	dt	<=	160	;
						10'd241	:	dt	<=	96	;
						10'd242	:	dt	<=	183	;
						10'd243	:	dt	<=	178	;
						10'd244	:	dt	<=	107	;
						10'd245	:	dt	<=	165	;
						10'd246	:	dt	<=	206	;
						10'd247	:	dt	<=	197	;
						10'd248	:	dt	<=	197	;
						10'd249	:	dt	<=	197	;
						10'd250	:	dt	<=	195	;
						10'd251	:	dt	<=	192	;
						10'd252	:	dt	<=	188	;
						10'd253	:	dt	<=	192	;
						10'd254	:	dt	<=	195	;
						10'd255	:	dt	<=	198	;
						10'd256	:	dt	<=	202	;
						10'd257	:	dt	<=	204	;
						10'd258	:	dt	<=	206	;
						10'd259	:	dt	<=	207	;
						10'd260	:	dt	<=	210	;
						10'd261	:	dt	<=	211	;
						10'd262	:	dt	<=	209	;
						10'd263	:	dt	<=	219	;
						10'd264	:	dt	<=	183	;
						10'd265	:	dt	<=	111	;
						10'd266	:	dt	<=	204	;
						10'd267	:	dt	<=	197	;
						10'd268	:	dt	<=	114	;
						10'd269	:	dt	<=	123	;
						10'd270	:	dt	<=	208	;
						10'd271	:	dt	<=	174	;
						10'd272	:	dt	<=	109	;
						10'd273	:	dt	<=	176	;
						10'd274	:	dt	<=	209	;
						10'd275	:	dt	<=	200	;
						10'd276	:	dt	<=	199	;
						10'd277	:	dt	<=	198	;
						10'd278	:	dt	<=	196	;
						10'd279	:	dt	<=	194	;
						10'd280	:	dt	<=	190	;
						10'd281	:	dt	<=	194	;
						10'd282	:	dt	<=	197	;
						10'd283	:	dt	<=	200	;
						10'd284	:	dt	<=	203	;
						10'd285	:	dt	<=	206	;
						10'd286	:	dt	<=	207	;
						10'd287	:	dt	<=	209	;
						10'd288	:	dt	<=	212	;
						10'd289	:	dt	<=	212	;
						10'd290	:	dt	<=	219	;
						10'd291	:	dt	<=	232	;
						10'd292	:	dt	<=	195	;
						10'd293	:	dt	<=	146	;
						10'd294	:	dt	<=	151	;
						10'd295	:	dt	<=	115	;
						10'd296	:	dt	<=	72	;
						10'd297	:	dt	<=	144	;
						10'd298	:	dt	<=	193	;
						10'd299	:	dt	<=	158	;
						10'd300	:	dt	<=	102	;
						10'd301	:	dt	<=	188	;
						10'd302	:	dt	<=	208	;
						10'd303	:	dt	<=	200	;
						10'd304	:	dt	<=	199	;
						10'd305	:	dt	<=	199	;
						10'd306	:	dt	<=	197	;
						10'd307	:	dt	<=	196	;
						10'd308	:	dt	<=	191	;
						10'd309	:	dt	<=	195	;
						10'd310	:	dt	<=	197	;
						10'd311	:	dt	<=	202	;
						10'd312	:	dt	<=	205	;
						10'd313	:	dt	<=	207	;
						10'd314	:	dt	<=	211	;
						10'd315	:	dt	<=	211	;
						10'd316	:	dt	<=	213	;
						10'd317	:	dt	<=	210	;
						10'd318	:	dt	<=	181	;
						10'd319	:	dt	<=	202	;
						10'd320	:	dt	<=	217	;
						10'd321	:	dt	<=	182	;
						10'd322	:	dt	<=	129	;
						10'd323	:	dt	<=	102	;
						10'd324	:	dt	<=	85	;
						10'd325	:	dt	<=	139	;
						10'd326	:	dt	<=	154	;
						10'd327	:	dt	<=	123	;
						10'd328	:	dt	<=	103	;
						10'd329	:	dt	<=	205	;
						10'd330	:	dt	<=	204	;
						10'd331	:	dt	<=	203	;
						10'd332	:	dt	<=	203	;
						10'd333	:	dt	<=	202	;
						10'd334	:	dt	<=	200	;
						10'd335	:	dt	<=	198	;
						10'd336	:	dt	<=	193	;
						10'd337	:	dt	<=	196	;
						10'd338	:	dt	<=	200	;
						10'd339	:	dt	<=	204	;
						10'd340	:	dt	<=	207	;
						10'd341	:	dt	<=	209	;
						10'd342	:	dt	<=	212	;
						10'd343	:	dt	<=	211	;
						10'd344	:	dt	<=	227	;
						10'd345	:	dt	<=	221	;
						10'd346	:	dt	<=	152	;
						10'd347	:	dt	<=	154	;
						10'd348	:	dt	<=	223	;
						10'd349	:	dt	<=	171	;
						10'd350	:	dt	<=	159	;
						10'd351	:	dt	<=	151	;
						10'd352	:	dt	<=	143	;
						10'd353	:	dt	<=	149	;
						10'd354	:	dt	<=	116	;
						10'd355	:	dt	<=	97	;
						10'd356	:	dt	<=	134	;
						10'd357	:	dt	<=	218	;
						10'd358	:	dt	<=	204	;
						10'd359	:	dt	<=	205	;
						10'd360	:	dt	<=	204	;
						10'd361	:	dt	<=	203	;
						10'd362	:	dt	<=	201	;
						10'd363	:	dt	<=	199	;
						10'd364	:	dt	<=	193	;
						10'd365	:	dt	<=	197	;
						10'd366	:	dt	<=	203	;
						10'd367	:	dt	<=	205	;
						10'd368	:	dt	<=	208	;
						10'd369	:	dt	<=	211	;
						10'd370	:	dt	<=	211	;
						10'd371	:	dt	<=	219	;
						10'd372	:	dt	<=	243	;
						10'd373	:	dt	<=	232	;
						10'd374	:	dt	<=	176	;
						10'd375	:	dt	<=	159	;
						10'd376	:	dt	<=	192	;
						10'd377	:	dt	<=	183	;
						10'd378	:	dt	<=	178	;
						10'd379	:	dt	<=	163	;
						10'd380	:	dt	<=	174	;
						10'd381	:	dt	<=	160	;
						10'd382	:	dt	<=	95	;
						10'd383	:	dt	<=	77	;
						10'd384	:	dt	<=	172	;
						10'd385	:	dt	<=	217	;
						10'd386	:	dt	<=	206	;
						10'd387	:	dt	<=	206	;
						10'd388	:	dt	<=	205	;
						10'd389	:	dt	<=	204	;
						10'd390	:	dt	<=	202	;
						10'd391	:	dt	<=	200	;
						10'd392	:	dt	<=	196	;
						10'd393	:	dt	<=	199	;
						10'd394	:	dt	<=	204	;
						10'd395	:	dt	<=	206	;
						10'd396	:	dt	<=	210	;
						10'd397	:	dt	<=	213	;
						10'd398	:	dt	<=	210	;
						10'd399	:	dt	<=	233	;
						10'd400	:	dt	<=	228	;
						10'd401	:	dt	<=	236	;
						10'd402	:	dt	<=	177	;
						10'd403	:	dt	<=	149	;
						10'd404	:	dt	<=	209	;
						10'd405	:	dt	<=	193	;
						10'd406	:	dt	<=	159	;
						10'd407	:	dt	<=	158	;
						10'd408	:	dt	<=	160	;
						10'd409	:	dt	<=	139	;
						10'd410	:	dt	<=	110	;
						10'd411	:	dt	<=	70	;
						10'd412	:	dt	<=	181	;
						10'd413	:	dt	<=	218	;
						10'd414	:	dt	<=	208	;
						10'd415	:	dt	<=	208	;
						10'd416	:	dt	<=	206	;
						10'd417	:	dt	<=	204	;
						10'd418	:	dt	<=	204	;
						10'd419	:	dt	<=	203	;
						10'd420	:	dt	<=	197	;
						10'd421	:	dt	<=	200	;
						10'd422	:	dt	<=	205	;
						10'd423	:	dt	<=	208	;
						10'd424	:	dt	<=	210	;
						10'd425	:	dt	<=	213	;
						10'd426	:	dt	<=	213	;
						10'd427	:	dt	<=	248	;
						10'd428	:	dt	<=	221	;
						10'd429	:	dt	<=	208	;
						10'd430	:	dt	<=	192	;
						10'd431	:	dt	<=	126	;
						10'd432	:	dt	<=	175	;
						10'd433	:	dt	<=	164	;
						10'd434	:	dt	<=	87	;
						10'd435	:	dt	<=	91	;
						10'd436	:	dt	<=	159	;
						10'd437	:	dt	<=	151	;
						10'd438	:	dt	<=	131	;
						10'd439	:	dt	<=	77	;
						10'd440	:	dt	<=	175	;
						10'd441	:	dt	<=	221	;
						10'd442	:	dt	<=	209	;
						10'd443	:	dt	<=	209	;
						10'd444	:	dt	<=	207	;
						10'd445	:	dt	<=	205	;
						10'd446	:	dt	<=	206	;
						10'd447	:	dt	<=	203	;
						10'd448	:	dt	<=	198	;
						10'd449	:	dt	<=	202	;
						10'd450	:	dt	<=	206	;
						10'd451	:	dt	<=	210	;
						10'd452	:	dt	<=	213	;
						10'd453	:	dt	<=	213	;
						10'd454	:	dt	<=	222	;
						10'd455	:	dt	<=	241	;
						10'd456	:	dt	<=	201	;
						10'd457	:	dt	<=	192	;
						10'd458	:	dt	<=	193	;
						10'd459	:	dt	<=	104	;
						10'd460	:	dt	<=	76	;
						10'd461	:	dt	<=	79	;
						10'd462	:	dt	<=	56	;
						10'd463	:	dt	<=	55	;
						10'd464	:	dt	<=	155	;
						10'd465	:	dt	<=	189	;
						10'd466	:	dt	<=	145	;
						10'd467	:	dt	<=	95	;
						10'd468	:	dt	<=	117	;
						10'd469	:	dt	<=	221	;
						10'd470	:	dt	<=	210	;
						10'd471	:	dt	<=	210	;
						10'd472	:	dt	<=	209	;
						10'd473	:	dt	<=	208	;
						10'd474	:	dt	<=	205	;
						10'd475	:	dt	<=	204	;
						10'd476	:	dt	<=	199	;
						10'd477	:	dt	<=	203	;
						10'd478	:	dt	<=	206	;
						10'd479	:	dt	<=	210	;
						10'd480	:	dt	<=	214	;
						10'd481	:	dt	<=	216	;
						10'd482	:	dt	<=	220	;
						10'd483	:	dt	<=	252	;
						10'd484	:	dt	<=	236	;
						10'd485	:	dt	<=	214	;
						10'd486	:	dt	<=	177	;
						10'd487	:	dt	<=	147	;
						10'd488	:	dt	<=	100	;
						10'd489	:	dt	<=	56	;
						10'd490	:	dt	<=	100	;
						10'd491	:	dt	<=	177	;
						10'd492	:	dt	<=	189	;
						10'd493	:	dt	<=	198	;
						10'd494	:	dt	<=	163	;
						10'd495	:	dt	<=	115	;
						10'd496	:	dt	<=	75	;
						10'd497	:	dt	<=	185	;
						10'd498	:	dt	<=	219	;
						10'd499	:	dt	<=	210	;
						10'd500	:	dt	<=	211	;
						10'd501	:	dt	<=	209	;
						10'd502	:	dt	<=	207	;
						10'd503	:	dt	<=	205	;
						10'd504	:	dt	<=	199	;
						10'd505	:	dt	<=	204	;
						10'd506	:	dt	<=	208	;
						10'd507	:	dt	<=	211	;
						10'd508	:	dt	<=	214	;
						10'd509	:	dt	<=	215	;
						10'd510	:	dt	<=	223	;
						10'd511	:	dt	<=	254	;
						10'd512	:	dt	<=	243	;
						10'd513	:	dt	<=	211	;
						10'd514	:	dt	<=	170	;
						10'd515	:	dt	<=	188	;
						10'd516	:	dt	<=	120	;
						10'd517	:	dt	<=	88	;
						10'd518	:	dt	<=	199	;
						10'd519	:	dt	<=	233	;
						10'd520	:	dt	<=	211	;
						10'd521	:	dt	<=	180	;
						10'd522	:	dt	<=	158	;
						10'd523	:	dt	<=	118	;
						10'd524	:	dt	<=	83	;
						10'd525	:	dt	<=	172	;
						10'd526	:	dt	<=	223	;
						10'd527	:	dt	<=	211	;
						10'd528	:	dt	<=	211	;
						10'd529	:	dt	<=	211	;
						10'd530	:	dt	<=	209	;
						10'd531	:	dt	<=	205	;
						10'd532	:	dt	<=	200	;
						10'd533	:	dt	<=	206	;
						10'd534	:	dt	<=	210	;
						10'd535	:	dt	<=	212	;
						10'd536	:	dt	<=	215	;
						10'd537	:	dt	<=	217	;
						10'd538	:	dt	<=	224	;
						10'd539	:	dt	<=	254	;
						10'd540	:	dt	<=	246	;
						10'd541	:	dt	<=	202	;
						10'd542	:	dt	<=	167	;
						10'd543	:	dt	<=	153	;
						10'd544	:	dt	<=	104	;
						10'd545	:	dt	<=	159	;
						10'd546	:	dt	<=	236	;
						10'd547	:	dt	<=	211	;
						10'd548	:	dt	<=	186	;
						10'd549	:	dt	<=	172	;
						10'd550	:	dt	<=	125	;
						10'd551	:	dt	<=	116	;
						10'd552	:	dt	<=	86	;
						10'd553	:	dt	<=	197	;
						10'd554	:	dt	<=	219	;
						10'd555	:	dt	<=	213	;
						10'd556	:	dt	<=	213	;
						10'd557	:	dt	<=	211	;
						10'd558	:	dt	<=	209	;
						10'd559	:	dt	<=	206	;
						10'd560	:	dt	<=	202	;
						10'd561	:	dt	<=	206	;
						10'd562	:	dt	<=	211	;
						10'd563	:	dt	<=	213	;
						10'd564	:	dt	<=	216	;
						10'd565	:	dt	<=	218	;
						10'd566	:	dt	<=	224	;
						10'd567	:	dt	<=	252	;
						10'd568	:	dt	<=	240	;
						10'd569	:	dt	<=	202	;
						10'd570	:	dt	<=	197	;
						10'd571	:	dt	<=	141	;
						10'd572	:	dt	<=	159	;
						10'd573	:	dt	<=	242	;
						10'd574	:	dt	<=	222	;
						10'd575	:	dt	<=	185	;
						10'd576	:	dt	<=	158	;
						10'd577	:	dt	<=	171	;
						10'd578	:	dt	<=	121	;
						10'd579	:	dt	<=	91	;
						10'd580	:	dt	<=	102	;
						10'd581	:	dt	<=	223	;
						10'd582	:	dt	<=	215	;
						10'd583	:	dt	<=	215	;
						10'd584	:	dt	<=	214	;
						10'd585	:	dt	<=	213	;
						10'd586	:	dt	<=	210	;
						10'd587	:	dt	<=	209	;
						10'd588	:	dt	<=	203	;
						10'd589	:	dt	<=	207	;
						10'd590	:	dt	<=	212	;
						10'd591	:	dt	<=	215	;
						10'd592	:	dt	<=	219	;
						10'd593	:	dt	<=	220	;
						10'd594	:	dt	<=	224	;
						10'd595	:	dt	<=	248	;
						10'd596	:	dt	<=	238	;
						10'd597	:	dt	<=	212	;
						10'd598	:	dt	<=	204	;
						10'd599	:	dt	<=	149	;
						10'd600	:	dt	<=	201	;
						10'd601	:	dt	<=	241	;
						10'd602	:	dt	<=	207	;
						10'd603	:	dt	<=	185	;
						10'd604	:	dt	<=	166	;
						10'd605	:	dt	<=	162	;
						10'd606	:	dt	<=	139	;
						10'd607	:	dt	<=	69	;
						10'd608	:	dt	<=	143	;
						10'd609	:	dt	<=	231	;
						10'd610	:	dt	<=	216	;
						10'd611	:	dt	<=	216	;
						10'd612	:	dt	<=	216	;
						10'd613	:	dt	<=	213	;
						10'd614	:	dt	<=	212	;
						10'd615	:	dt	<=	209	;
						10'd616	:	dt	<=	203	;
						10'd617	:	dt	<=	208	;
						10'd618	:	dt	<=	212	;
						10'd619	:	dt	<=	216	;
						10'd620	:	dt	<=	219	;
						10'd621	:	dt	<=	221	;
						10'd622	:	dt	<=	224	;
						10'd623	:	dt	<=	238	;
						10'd624	:	dt	<=	233	;
						10'd625	:	dt	<=	214	;
						10'd626	:	dt	<=	204	;
						10'd627	:	dt	<=	155	;
						10'd628	:	dt	<=	191	;
						10'd629	:	dt	<=	217	;
						10'd630	:	dt	<=	193	;
						10'd631	:	dt	<=	180	;
						10'd632	:	dt	<=	155	;
						10'd633	:	dt	<=	141	;
						10'd634	:	dt	<=	120	;
						10'd635	:	dt	<=	71	;
						10'd636	:	dt	<=	200	;
						10'd637	:	dt	<=	224	;
						10'd638	:	dt	<=	217	;
						10'd639	:	dt	<=	218	;
						10'd640	:	dt	<=	216	;
						10'd641	:	dt	<=	214	;
						10'd642	:	dt	<=	212	;
						10'd643	:	dt	<=	210	;
						10'd644	:	dt	<=	204	;
						10'd645	:	dt	<=	209	;
						10'd646	:	dt	<=	213	;
						10'd647	:	dt	<=	217	;
						10'd648	:	dt	<=	217	;
						10'd649	:	dt	<=	223	;
						10'd650	:	dt	<=	227	;
						10'd651	:	dt	<=	237	;
						10'd652	:	dt	<=	232	;
						10'd653	:	dt	<=	216	;
						10'd654	:	dt	<=	196	;
						10'd655	:	dt	<=	157	;
						10'd656	:	dt	<=	155	;
						10'd657	:	dt	<=	181	;
						10'd658	:	dt	<=	170	;
						10'd659	:	dt	<=	153	;
						10'd660	:	dt	<=	131	;
						10'd661	:	dt	<=	125	;
						10'd662	:	dt	<=	76	;
						10'd663	:	dt	<=	133	;
						10'd664	:	dt	<=	233	;
						10'd665	:	dt	<=	218	;
						10'd666	:	dt	<=	220	;
						10'd667	:	dt	<=	219	;
						10'd668	:	dt	<=	217	;
						10'd669	:	dt	<=	215	;
						10'd670	:	dt	<=	213	;
						10'd671	:	dt	<=	211	;
						10'd672	:	dt	<=	203	;
						10'd673	:	dt	<=	207	;
						10'd674	:	dt	<=	212	;
						10'd675	:	dt	<=	214	;
						10'd676	:	dt	<=	226	;
						10'd677	:	dt	<=	201	;
						10'd678	:	dt	<=	96	;
						10'd679	:	dt	<=	184	;
						10'd680	:	dt	<=	228	;
						10'd681	:	dt	<=	212	;
						10'd682	:	dt	<=	163	;
						10'd683	:	dt	<=	128	;
						10'd684	:	dt	<=	131	;
						10'd685	:	dt	<=	144	;
						10'd686	:	dt	<=	163	;
						10'd687	:	dt	<=	141	;
						10'd688	:	dt	<=	117	;
						10'd689	:	dt	<=	82	;
						10'd690	:	dt	<=	82	;
						10'd691	:	dt	<=	218	;
						10'd692	:	dt	<=	225	;
						10'd693	:	dt	<=	221	;
						10'd694	:	dt	<=	220	;
						10'd695	:	dt	<=	219	;
						10'd696	:	dt	<=	218	;
						10'd697	:	dt	<=	216	;
						10'd698	:	dt	<=	213	;
						10'd699	:	dt	<=	211	;
						10'd700	:	dt	<=	202	;
						10'd701	:	dt	<=	205	;
						10'd702	:	dt	<=	209	;
						10'd703	:	dt	<=	219	;
						10'd704	:	dt	<=	212	;
						10'd705	:	dt	<=	104	;
						10'd706	:	dt	<=	61	;
						10'd707	:	dt	<=	76	;
						10'd708	:	dt	<=	163	;
						10'd709	:	dt	<=	179	;
						10'd710	:	dt	<=	140	;
						10'd711	:	dt	<=	133	;
						10'd712	:	dt	<=	141	;
						10'd713	:	dt	<=	145	;
						10'd714	:	dt	<=	168	;
						10'd715	:	dt	<=	133	;
						10'd716	:	dt	<=	98	;
						10'd717	:	dt	<=	67	;
						10'd718	:	dt	<=	183	;
						10'd719	:	dt	<=	231	;
						10'd720	:	dt	<=	219	;
						10'd721	:	dt	<=	221	;
						10'd722	:	dt	<=	220	;
						10'd723	:	dt	<=	219	;
						10'd724	:	dt	<=	217	;
						10'd725	:	dt	<=	214	;
						10'd726	:	dt	<=	212	;
						10'd727	:	dt	<=	210	;
						10'd728	:	dt	<=	203	;
						10'd729	:	dt	<=	207	;
						10'd730	:	dt	<=	213	;
						10'd731	:	dt	<=	217	;
						10'd732	:	dt	<=	114	;
						10'd733	:	dt	<=	65	;
						10'd734	:	dt	<=	79	;
						10'd735	:	dt	<=	67	;
						10'd736	:	dt	<=	76	;
						10'd737	:	dt	<=	138	;
						10'd738	:	dt	<=	157	;
						10'd739	:	dt	<=	150	;
						10'd740	:	dt	<=	144	;
						10'd741	:	dt	<=	145	;
						10'd742	:	dt	<=	154	;
						10'd743	:	dt	<=	118	;
						10'd744	:	dt	<=	68	;
						10'd745	:	dt	<=	150	;
						10'd746	:	dt	<=	237	;
						10'd747	:	dt	<=	221	;
						10'd748	:	dt	<=	222	;
						10'd749	:	dt	<=	221	;
						10'd750	:	dt	<=	220	;
						10'd751	:	dt	<=	218	;
						10'd752	:	dt	<=	217	;
						10'd753	:	dt	<=	214	;
						10'd754	:	dt	<=	213	;
						10'd755	:	dt	<=	210	;
						10'd756	:	dt	<=	203	;
						10'd757	:	dt	<=	206	;
						10'd758	:	dt	<=	221	;
						10'd759	:	dt	<=	137	;
						10'd760	:	dt	<=	72	;
						10'd761	:	dt	<=	82	;
						10'd762	:	dt	<=	66	;
						10'd763	:	dt	<=	71	;
						10'd764	:	dt	<=	65	;
						10'd765	:	dt	<=	72	;
						10'd766	:	dt	<=	118	;
						10'd767	:	dt	<=	129	;
						10'd768	:	dt	<=	133	;
						10'd769	:	dt	<=	131	;
						10'd770	:	dt	<=	119	;
						10'd771	:	dt	<=	89	;
						10'd772	:	dt	<=	91	;
						10'd773	:	dt	<=	223	;
						10'd774	:	dt	<=	227	;
						10'd775	:	dt	<=	224	;
						10'd776	:	dt	<=	223	;
						10'd777	:	dt	<=	221	;
						10'd778	:	dt	<=	220	;
						10'd779	:	dt	<=	219	;
						10'd780	:	dt	<=	218	;
						10'd781	:	dt	<=	216	;
						10'd782	:	dt	<=	214	;
						10'd783	:	dt	<=	212	;
					endcase
				end
				5'd21	:	begin
					case (cnt)
						10'd0	:	dt	<=	72	;
						10'd1	:	dt	<=	79	;
						10'd2	:	dt	<=	87	;
						10'd3	:	dt	<=	101	;
						10'd4	:	dt	<=	115	;
						10'd5	:	dt	<=	124	;
						10'd6	:	dt	<=	131	;
						10'd7	:	dt	<=	135	;
						10'd8	:	dt	<=	139	;
						10'd9	:	dt	<=	142	;
						10'd10	:	dt	<=	144	;
						10'd11	:	dt	<=	147	;
						10'd12	:	dt	<=	150	;
						10'd13	:	dt	<=	153	;
						10'd14	:	dt	<=	156	;
						10'd15	:	dt	<=	159	;
						10'd16	:	dt	<=	160	;
						10'd17	:	dt	<=	162	;
						10'd18	:	dt	<=	164	;
						10'd19	:	dt	<=	165	;
						10'd20	:	dt	<=	166	;
						10'd21	:	dt	<=	166	;
						10'd22	:	dt	<=	167	;
						10'd23	:	dt	<=	167	;
						10'd24	:	dt	<=	168	;
						10'd25	:	dt	<=	168	;
						10'd26	:	dt	<=	168	;
						10'd27	:	dt	<=	167	;
						10'd28	:	dt	<=	73	;
						10'd29	:	dt	<=	80	;
						10'd30	:	dt	<=	89	;
						10'd31	:	dt	<=	104	;
						10'd32	:	dt	<=	117	;
						10'd33	:	dt	<=	126	;
						10'd34	:	dt	<=	132	;
						10'd35	:	dt	<=	136	;
						10'd36	:	dt	<=	140	;
						10'd37	:	dt	<=	143	;
						10'd38	:	dt	<=	146	;
						10'd39	:	dt	<=	149	;
						10'd40	:	dt	<=	152	;
						10'd41	:	dt	<=	155	;
						10'd42	:	dt	<=	150	;
						10'd43	:	dt	<=	160	;
						10'd44	:	dt	<=	163	;
						10'd45	:	dt	<=	164	;
						10'd46	:	dt	<=	165	;
						10'd47	:	dt	<=	166	;
						10'd48	:	dt	<=	168	;
						10'd49	:	dt	<=	169	;
						10'd50	:	dt	<=	169	;
						10'd51	:	dt	<=	169	;
						10'd52	:	dt	<=	170	;
						10'd53	:	dt	<=	169	;
						10'd54	:	dt	<=	169	;
						10'd55	:	dt	<=	169	;
						10'd56	:	dt	<=	75	;
						10'd57	:	dt	<=	82	;
						10'd58	:	dt	<=	90	;
						10'd59	:	dt	<=	107	;
						10'd60	:	dt	<=	119	;
						10'd61	:	dt	<=	128	;
						10'd62	:	dt	<=	134	;
						10'd63	:	dt	<=	138	;
						10'd64	:	dt	<=	142	;
						10'd65	:	dt	<=	145	;
						10'd66	:	dt	<=	147	;
						10'd67	:	dt	<=	152	;
						10'd68	:	dt	<=	159	;
						10'd69	:	dt	<=	162	;
						10'd70	:	dt	<=	105	;
						10'd71	:	dt	<=	153	;
						10'd72	:	dt	<=	165	;
						10'd73	:	dt	<=	167	;
						10'd74	:	dt	<=	168	;
						10'd75	:	dt	<=	168	;
						10'd76	:	dt	<=	170	;
						10'd77	:	dt	<=	171	;
						10'd78	:	dt	<=	171	;
						10'd79	:	dt	<=	171	;
						10'd80	:	dt	<=	171	;
						10'd81	:	dt	<=	172	;
						10'd82	:	dt	<=	171	;
						10'd83	:	dt	<=	171	;
						10'd84	:	dt	<=	76	;
						10'd85	:	dt	<=	84	;
						10'd86	:	dt	<=	92	;
						10'd87	:	dt	<=	109	;
						10'd88	:	dt	<=	121	;
						10'd89	:	dt	<=	128	;
						10'd90	:	dt	<=	135	;
						10'd91	:	dt	<=	140	;
						10'd92	:	dt	<=	143	;
						10'd93	:	dt	<=	146	;
						10'd94	:	dt	<=	150	;
						10'd95	:	dt	<=	153	;
						10'd96	:	dt	<=	167	;
						10'd97	:	dt	<=	160	;
						10'd98	:	dt	<=	101	;
						10'd99	:	dt	<=	149	;
						10'd100	:	dt	<=	168	;
						10'd101	:	dt	<=	168	;
						10'd102	:	dt	<=	169	;
						10'd103	:	dt	<=	171	;
						10'd104	:	dt	<=	173	;
						10'd105	:	dt	<=	173	;
						10'd106	:	dt	<=	172	;
						10'd107	:	dt	<=	172	;
						10'd108	:	dt	<=	173	;
						10'd109	:	dt	<=	173	;
						10'd110	:	dt	<=	173	;
						10'd111	:	dt	<=	173	;
						10'd112	:	dt	<=	77	;
						10'd113	:	dt	<=	85	;
						10'd114	:	dt	<=	94	;
						10'd115	:	dt	<=	111	;
						10'd116	:	dt	<=	122	;
						10'd117	:	dt	<=	130	;
						10'd118	:	dt	<=	136	;
						10'd119	:	dt	<=	141	;
						10'd120	:	dt	<=	146	;
						10'd121	:	dt	<=	149	;
						10'd122	:	dt	<=	152	;
						10'd123	:	dt	<=	155	;
						10'd124	:	dt	<=	170	;
						10'd125	:	dt	<=	159	;
						10'd126	:	dt	<=	106	;
						10'd127	:	dt	<=	145	;
						10'd128	:	dt	<=	168	;
						10'd129	:	dt	<=	171	;
						10'd130	:	dt	<=	171	;
						10'd131	:	dt	<=	172	;
						10'd132	:	dt	<=	175	;
						10'd133	:	dt	<=	175	;
						10'd134	:	dt	<=	175	;
						10'd135	:	dt	<=	175	;
						10'd136	:	dt	<=	177	;
						10'd137	:	dt	<=	175	;
						10'd138	:	dt	<=	175	;
						10'd139	:	dt	<=	174	;
						10'd140	:	dt	<=	78	;
						10'd141	:	dt	<=	86	;
						10'd142	:	dt	<=	96	;
						10'd143	:	dt	<=	112	;
						10'd144	:	dt	<=	123	;
						10'd145	:	dt	<=	132	;
						10'd146	:	dt	<=	137	;
						10'd147	:	dt	<=	141	;
						10'd148	:	dt	<=	146	;
						10'd149	:	dt	<=	150	;
						10'd150	:	dt	<=	152	;
						10'd151	:	dt	<=	156	;
						10'd152	:	dt	<=	173	;
						10'd153	:	dt	<=	165	;
						10'd154	:	dt	<=	112	;
						10'd155	:	dt	<=	143	;
						10'd156	:	dt	<=	170	;
						10'd157	:	dt	<=	171	;
						10'd158	:	dt	<=	173	;
						10'd159	:	dt	<=	173	;
						10'd160	:	dt	<=	177	;
						10'd161	:	dt	<=	177	;
						10'd162	:	dt	<=	171	;
						10'd163	:	dt	<=	161	;
						10'd164	:	dt	<=	176	;
						10'd165	:	dt	<=	177	;
						10'd166	:	dt	<=	177	;
						10'd167	:	dt	<=	177	;
						10'd168	:	dt	<=	79	;
						10'd169	:	dt	<=	88	;
						10'd170	:	dt	<=	98	;
						10'd171	:	dt	<=	115	;
						10'd172	:	dt	<=	124	;
						10'd173	:	dt	<=	133	;
						10'd174	:	dt	<=	139	;
						10'd175	:	dt	<=	144	;
						10'd176	:	dt	<=	148	;
						10'd177	:	dt	<=	150	;
						10'd178	:	dt	<=	153	;
						10'd179	:	dt	<=	157	;
						10'd180	:	dt	<=	175	;
						10'd181	:	dt	<=	165	;
						10'd182	:	dt	<=	117	;
						10'd183	:	dt	<=	136	;
						10'd184	:	dt	<=	172	;
						10'd185	:	dt	<=	174	;
						10'd186	:	dt	<=	176	;
						10'd187	:	dt	<=	176	;
						10'd188	:	dt	<=	177	;
						10'd189	:	dt	<=	175	;
						10'd190	:	dt	<=	145	;
						10'd191	:	dt	<=	108	;
						10'd192	:	dt	<=	164	;
						10'd193	:	dt	<=	179	;
						10'd194	:	dt	<=	179	;
						10'd195	:	dt	<=	179	;
						10'd196	:	dt	<=	81	;
						10'd197	:	dt	<=	89	;
						10'd198	:	dt	<=	100	;
						10'd199	:	dt	<=	117	;
						10'd200	:	dt	<=	126	;
						10'd201	:	dt	<=	135	;
						10'd202	:	dt	<=	140	;
						10'd203	:	dt	<=	145	;
						10'd204	:	dt	<=	149	;
						10'd205	:	dt	<=	150	;
						10'd206	:	dt	<=	154	;
						10'd207	:	dt	<=	158	;
						10'd208	:	dt	<=	176	;
						10'd209	:	dt	<=	165	;
						10'd210	:	dt	<=	120	;
						10'd211	:	dt	<=	124	;
						10'd212	:	dt	<=	173	;
						10'd213	:	dt	<=	174	;
						10'd214	:	dt	<=	177	;
						10'd215	:	dt	<=	177	;
						10'd216	:	dt	<=	179	;
						10'd217	:	dt	<=	163	;
						10'd218	:	dt	<=	126	;
						10'd219	:	dt	<=	110	;
						10'd220	:	dt	<=	175	;
						10'd221	:	dt	<=	181	;
						10'd222	:	dt	<=	180	;
						10'd223	:	dt	<=	180	;
						10'd224	:	dt	<=	83	;
						10'd225	:	dt	<=	90	;
						10'd226	:	dt	<=	101	;
						10'd227	:	dt	<=	118	;
						10'd228	:	dt	<=	126	;
						10'd229	:	dt	<=	134	;
						10'd230	:	dt	<=	141	;
						10'd231	:	dt	<=	147	;
						10'd232	:	dt	<=	150	;
						10'd233	:	dt	<=	151	;
						10'd234	:	dt	<=	155	;
						10'd235	:	dt	<=	160	;
						10'd236	:	dt	<=	181	;
						10'd237	:	dt	<=	167	;
						10'd238	:	dt	<=	121	;
						10'd239	:	dt	<=	121	;
						10'd240	:	dt	<=	174	;
						10'd241	:	dt	<=	175	;
						10'd242	:	dt	<=	178	;
						10'd243	:	dt	<=	180	;
						10'd244	:	dt	<=	177	;
						10'd245	:	dt	<=	144	;
						10'd246	:	dt	<=	108	;
						10'd247	:	dt	<=	155	;
						10'd248	:	dt	<=	183	;
						10'd249	:	dt	<=	182	;
						10'd250	:	dt	<=	182	;
						10'd251	:	dt	<=	181	;
						10'd252	:	dt	<=	84	;
						10'd253	:	dt	<=	91	;
						10'd254	:	dt	<=	104	;
						10'd255	:	dt	<=	120	;
						10'd256	:	dt	<=	129	;
						10'd257	:	dt	<=	137	;
						10'd258	:	dt	<=	142	;
						10'd259	:	dt	<=	148	;
						10'd260	:	dt	<=	151	;
						10'd261	:	dt	<=	152	;
						10'd262	:	dt	<=	157	;
						10'd263	:	dt	<=	160	;
						10'd264	:	dt	<=	188	;
						10'd265	:	dt	<=	170	;
						10'd266	:	dt	<=	127	;
						10'd267	:	dt	<=	126	;
						10'd268	:	dt	<=	175	;
						10'd269	:	dt	<=	176	;
						10'd270	:	dt	<=	179	;
						10'd271	:	dt	<=	176	;
						10'd272	:	dt	<=	156	;
						10'd273	:	dt	<=	124	;
						10'd274	:	dt	<=	127	;
						10'd275	:	dt	<=	181	;
						10'd276	:	dt	<=	184	;
						10'd277	:	dt	<=	183	;
						10'd278	:	dt	<=	183	;
						10'd279	:	dt	<=	182	;
						10'd280	:	dt	<=	84	;
						10'd281	:	dt	<=	92	;
						10'd282	:	dt	<=	107	;
						10'd283	:	dt	<=	121	;
						10'd284	:	dt	<=	130	;
						10'd285	:	dt	<=	138	;
						10'd286	:	dt	<=	143	;
						10'd287	:	dt	<=	148	;
						10'd288	:	dt	<=	151	;
						10'd289	:	dt	<=	154	;
						10'd290	:	dt	<=	162	;
						10'd291	:	dt	<=	147	;
						10'd292	:	dt	<=	172	;
						10'd293	:	dt	<=	152	;
						10'd294	:	dt	<=	121	;
						10'd295	:	dt	<=	122	;
						10'd296	:	dt	<=	176	;
						10'd297	:	dt	<=	177	;
						10'd298	:	dt	<=	181	;
						10'd299	:	dt	<=	171	;
						10'd300	:	dt	<=	137	;
						10'd301	:	dt	<=	107	;
						10'd302	:	dt	<=	170	;
						10'd303	:	dt	<=	184	;
						10'd304	:	dt	<=	185	;
						10'd305	:	dt	<=	185	;
						10'd306	:	dt	<=	185	;
						10'd307	:	dt	<=	184	;
						10'd308	:	dt	<=	86	;
						10'd309	:	dt	<=	93	;
						10'd310	:	dt	<=	108	;
						10'd311	:	dt	<=	121	;
						10'd312	:	dt	<=	131	;
						10'd313	:	dt	<=	138	;
						10'd314	:	dt	<=	144	;
						10'd315	:	dt	<=	149	;
						10'd316	:	dt	<=	152	;
						10'd317	:	dt	<=	161	;
						10'd318	:	dt	<=	159	;
						10'd319	:	dt	<=	128	;
						10'd320	:	dt	<=	121	;
						10'd321	:	dt	<=	112	;
						10'd322	:	dt	<=	107	;
						10'd323	:	dt	<=	122	;
						10'd324	:	dt	<=	177	;
						10'd325	:	dt	<=	178	;
						10'd326	:	dt	<=	179	;
						10'd327	:	dt	<=	159	;
						10'd328	:	dt	<=	115	;
						10'd329	:	dt	<=	139	;
						10'd330	:	dt	<=	185	;
						10'd331	:	dt	<=	185	;
						10'd332	:	dt	<=	186	;
						10'd333	:	dt	<=	186	;
						10'd334	:	dt	<=	185	;
						10'd335	:	dt	<=	185	;
						10'd336	:	dt	<=	87	;
						10'd337	:	dt	<=	95	;
						10'd338	:	dt	<=	110	;
						10'd339	:	dt	<=	122	;
						10'd340	:	dt	<=	131	;
						10'd341	:	dt	<=	139	;
						10'd342	:	dt	<=	145	;
						10'd343	:	dt	<=	151	;
						10'd344	:	dt	<=	162	;
						10'd345	:	dt	<=	177	;
						10'd346	:	dt	<=	136	;
						10'd347	:	dt	<=	121	;
						10'd348	:	dt	<=	91	;
						10'd349	:	dt	<=	84	;
						10'd350	:	dt	<=	92	;
						10'd351	:	dt	<=	122	;
						10'd352	:	dt	<=	161	;
						10'd353	:	dt	<=	165	;
						10'd354	:	dt	<=	162	;
						10'd355	:	dt	<=	128	;
						10'd356	:	dt	<=	109	;
						10'd357	:	dt	<=	178	;
						10'd358	:	dt	<=	186	;
						10'd359	:	dt	<=	187	;
						10'd360	:	dt	<=	187	;
						10'd361	:	dt	<=	187	;
						10'd362	:	dt	<=	186	;
						10'd363	:	dt	<=	186	;
						10'd364	:	dt	<=	88	;
						10'd365	:	dt	<=	95	;
						10'd366	:	dt	<=	111	;
						10'd367	:	dt	<=	123	;
						10'd368	:	dt	<=	132	;
						10'd369	:	dt	<=	139	;
						10'd370	:	dt	<=	146	;
						10'd371	:	dt	<=	152	;
						10'd372	:	dt	<=	186	;
						10'd373	:	dt	<=	189	;
						10'd374	:	dt	<=	166	;
						10'd375	:	dt	<=	139	;
						10'd376	:	dt	<=	93	;
						10'd377	:	dt	<=	72	;
						10'd378	:	dt	<=	85	;
						10'd379	:	dt	<=	112	;
						10'd380	:	dt	<=	141	;
						10'd381	:	dt	<=	143	;
						10'd382	:	dt	<=	126	;
						10'd383	:	dt	<=	97	;
						10'd384	:	dt	<=	154	;
						10'd385	:	dt	<=	186	;
						10'd386	:	dt	<=	186	;
						10'd387	:	dt	<=	187	;
						10'd388	:	dt	<=	187	;
						10'd389	:	dt	<=	188	;
						10'd390	:	dt	<=	187	;
						10'd391	:	dt	<=	186	;
						10'd392	:	dt	<=	88	;
						10'd393	:	dt	<=	96	;
						10'd394	:	dt	<=	113	;
						10'd395	:	dt	<=	124	;
						10'd396	:	dt	<=	132	;
						10'd397	:	dt	<=	140	;
						10'd398	:	dt	<=	146	;
						10'd399	:	dt	<=	158	;
						10'd400	:	dt	<=	192	;
						10'd401	:	dt	<=	197	;
						10'd402	:	dt	<=	195	;
						10'd403	:	dt	<=	140	;
						10'd404	:	dt	<=	95	;
						10'd405	:	dt	<=	73	;
						10'd406	:	dt	<=	80	;
						10'd407	:	dt	<=	100	;
						10'd408	:	dt	<=	118	;
						10'd409	:	dt	<=	120	;
						10'd410	:	dt	<=	99	;
						10'd411	:	dt	<=	116	;
						10'd412	:	dt	<=	183	;
						10'd413	:	dt	<=	188	;
						10'd414	:	dt	<=	188	;
						10'd415	:	dt	<=	188	;
						10'd416	:	dt	<=	188	;
						10'd417	:	dt	<=	189	;
						10'd418	:	dt	<=	189	;
						10'd419	:	dt	<=	189	;
						10'd420	:	dt	<=	89	;
						10'd421	:	dt	<=	97	;
						10'd422	:	dt	<=	114	;
						10'd423	:	dt	<=	124	;
						10'd424	:	dt	<=	133	;
						10'd425	:	dt	<=	140	;
						10'd426	:	dt	<=	147	;
						10'd427	:	dt	<=	167	;
						10'd428	:	dt	<=	174	;
						10'd429	:	dt	<=	163	;
						10'd430	:	dt	<=	170	;
						10'd431	:	dt	<=	128	;
						10'd432	:	dt	<=	93	;
						10'd433	:	dt	<=	79	;
						10'd434	:	dt	<=	77	;
						10'd435	:	dt	<=	91	;
						10'd436	:	dt	<=	102	;
						10'd437	:	dt	<=	103	;
						10'd438	:	dt	<=	92	;
						10'd439	:	dt	<=	170	;
						10'd440	:	dt	<=	188	;
						10'd441	:	dt	<=	189	;
						10'd442	:	dt	<=	188	;
						10'd443	:	dt	<=	189	;
						10'd444	:	dt	<=	189	;
						10'd445	:	dt	<=	189	;
						10'd446	:	dt	<=	190	;
						10'd447	:	dt	<=	189	;
						10'd448	:	dt	<=	90	;
						10'd449	:	dt	<=	98	;
						10'd450	:	dt	<=	115	;
						10'd451	:	dt	<=	125	;
						10'd452	:	dt	<=	133	;
						10'd453	:	dt	<=	141	;
						10'd454	:	dt	<=	147	;
						10'd455	:	dt	<=	184	;
						10'd456	:	dt	<=	165	;
						10'd457	:	dt	<=	121	;
						10'd458	:	dt	<=	138	;
						10'd459	:	dt	<=	136	;
						10'd460	:	dt	<=	104	;
						10'd461	:	dt	<=	83	;
						10'd462	:	dt	<=	78	;
						10'd463	:	dt	<=	82	;
						10'd464	:	dt	<=	89	;
						10'd465	:	dt	<=	84	;
						10'd466	:	dt	<=	118	;
						10'd467	:	dt	<=	187	;
						10'd468	:	dt	<=	188	;
						10'd469	:	dt	<=	189	;
						10'd470	:	dt	<=	190	;
						10'd471	:	dt	<=	190	;
						10'd472	:	dt	<=	190	;
						10'd473	:	dt	<=	190	;
						10'd474	:	dt	<=	190	;
						10'd475	:	dt	<=	189	;
						10'd476	:	dt	<=	91	;
						10'd477	:	dt	<=	99	;
						10'd478	:	dt	<=	116	;
						10'd479	:	dt	<=	125	;
						10'd480	:	dt	<=	134	;
						10'd481	:	dt	<=	142	;
						10'd482	:	dt	<=	151	;
						10'd483	:	dt	<=	183	;
						10'd484	:	dt	<=	140	;
						10'd485	:	dt	<=	113	;
						10'd486	:	dt	<=	117	;
						10'd487	:	dt	<=	151	;
						10'd488	:	dt	<=	116	;
						10'd489	:	dt	<=	90	;
						10'd490	:	dt	<=	80	;
						10'd491	:	dt	<=	76	;
						10'd492	:	dt	<=	81	;
						10'd493	:	dt	<=	80	;
						10'd494	:	dt	<=	145	;
						10'd495	:	dt	<=	188	;
						10'd496	:	dt	<=	189	;
						10'd497	:	dt	<=	190	;
						10'd498	:	dt	<=	190	;
						10'd499	:	dt	<=	190	;
						10'd500	:	dt	<=	190	;
						10'd501	:	dt	<=	191	;
						10'd502	:	dt	<=	192	;
						10'd503	:	dt	<=	190	;
						10'd504	:	dt	<=	91	;
						10'd505	:	dt	<=	101	;
						10'd506	:	dt	<=	118	;
						10'd507	:	dt	<=	125	;
						10'd508	:	dt	<=	135	;
						10'd509	:	dt	<=	141	;
						10'd510	:	dt	<=	162	;
						10'd511	:	dt	<=	183	;
						10'd512	:	dt	<=	153	;
						10'd513	:	dt	<=	142	;
						10'd514	:	dt	<=	138	;
						10'd515	:	dt	<=	172	;
						10'd516	:	dt	<=	131	;
						10'd517	:	dt	<=	110	;
						10'd518	:	dt	<=	89	;
						10'd519	:	dt	<=	77	;
						10'd520	:	dt	<=	76	;
						10'd521	:	dt	<=	79	;
						10'd522	:	dt	<=	154	;
						10'd523	:	dt	<=	189	;
						10'd524	:	dt	<=	191	;
						10'd525	:	dt	<=	192	;
						10'd526	:	dt	<=	191	;
						10'd527	:	dt	<=	191	;
						10'd528	:	dt	<=	191	;
						10'd529	:	dt	<=	191	;
						10'd530	:	dt	<=	192	;
						10'd531	:	dt	<=	190	;
						10'd532	:	dt	<=	91	;
						10'd533	:	dt	<=	102	;
						10'd534	:	dt	<=	117	;
						10'd535	:	dt	<=	125	;
						10'd536	:	dt	<=	135	;
						10'd537	:	dt	<=	143	;
						10'd538	:	dt	<=	174	;
						10'd539	:	dt	<=	183	;
						10'd540	:	dt	<=	166	;
						10'd541	:	dt	<=	141	;
						10'd542	:	dt	<=	174	;
						10'd543	:	dt	<=	194	;
						10'd544	:	dt	<=	139	;
						10'd545	:	dt	<=	124	;
						10'd546	:	dt	<=	94	;
						10'd547	:	dt	<=	76	;
						10'd548	:	dt	<=	76	;
						10'd549	:	dt	<=	81	;
						10'd550	:	dt	<=	168	;
						10'd551	:	dt	<=	189	;
						10'd552	:	dt	<=	191	;
						10'd553	:	dt	<=	192	;
						10'd554	:	dt	<=	193	;
						10'd555	:	dt	<=	193	;
						10'd556	:	dt	<=	193	;
						10'd557	:	dt	<=	193	;
						10'd558	:	dt	<=	192	;
						10'd559	:	dt	<=	191	;
						10'd560	:	dt	<=	92	;
						10'd561	:	dt	<=	103	;
						10'd562	:	dt	<=	119	;
						10'd563	:	dt	<=	126	;
						10'd564	:	dt	<=	136	;
						10'd565	:	dt	<=	143	;
						10'd566	:	dt	<=	184	;
						10'd567	:	dt	<=	193	;
						10'd568	:	dt	<=	164	;
						10'd569	:	dt	<=	147	;
						10'd570	:	dt	<=	205	;
						10'd571	:	dt	<=	178	;
						10'd572	:	dt	<=	135	;
						10'd573	:	dt	<=	120	;
						10'd574	:	dt	<=	94	;
						10'd575	:	dt	<=	76	;
						10'd576	:	dt	<=	75	;
						10'd577	:	dt	<=	85	;
						10'd578	:	dt	<=	180	;
						10'd579	:	dt	<=	191	;
						10'd580	:	dt	<=	192	;
						10'd581	:	dt	<=	192	;
						10'd582	:	dt	<=	193	;
						10'd583	:	dt	<=	193	;
						10'd584	:	dt	<=	193	;
						10'd585	:	dt	<=	193	;
						10'd586	:	dt	<=	193	;
						10'd587	:	dt	<=	192	;
						10'd588	:	dt	<=	93	;
						10'd589	:	dt	<=	104	;
						10'd590	:	dt	<=	119	;
						10'd591	:	dt	<=	127	;
						10'd592	:	dt	<=	136	;
						10'd593	:	dt	<=	143	;
						10'd594	:	dt	<=	190	;
						10'd595	:	dt	<=	184	;
						10'd596	:	dt	<=	157	;
						10'd597	:	dt	<=	157	;
						10'd598	:	dt	<=	197	;
						10'd599	:	dt	<=	163	;
						10'd600	:	dt	<=	130	;
						10'd601	:	dt	<=	113	;
						10'd602	:	dt	<=	100	;
						10'd603	:	dt	<=	79	;
						10'd604	:	dt	<=	75	;
						10'd605	:	dt	<=	104	;
						10'd606	:	dt	<=	189	;
						10'd607	:	dt	<=	192	;
						10'd608	:	dt	<=	192	;
						10'd609	:	dt	<=	192	;
						10'd610	:	dt	<=	193	;
						10'd611	:	dt	<=	193	;
						10'd612	:	dt	<=	194	;
						10'd613	:	dt	<=	194	;
						10'd614	:	dt	<=	193	;
						10'd615	:	dt	<=	193	;
						10'd616	:	dt	<=	92	;
						10'd617	:	dt	<=	104	;
						10'd618	:	dt	<=	118	;
						10'd619	:	dt	<=	127	;
						10'd620	:	dt	<=	137	;
						10'd621	:	dt	<=	144	;
						10'd622	:	dt	<=	183	;
						10'd623	:	dt	<=	170	;
						10'd624	:	dt	<=	166	;
						10'd625	:	dt	<=	158	;
						10'd626	:	dt	<=	193	;
						10'd627	:	dt	<=	158	;
						10'd628	:	dt	<=	144	;
						10'd629	:	dt	<=	110	;
						10'd630	:	dt	<=	91	;
						10'd631	:	dt	<=	79	;
						10'd632	:	dt	<=	75	;
						10'd633	:	dt	<=	138	;
						10'd634	:	dt	<=	190	;
						10'd635	:	dt	<=	192	;
						10'd636	:	dt	<=	192	;
						10'd637	:	dt	<=	192	;
						10'd638	:	dt	<=	193	;
						10'd639	:	dt	<=	194	;
						10'd640	:	dt	<=	195	;
						10'd641	:	dt	<=	194	;
						10'd642	:	dt	<=	193	;
						10'd643	:	dt	<=	194	;
						10'd644	:	dt	<=	92	;
						10'd645	:	dt	<=	106	;
						10'd646	:	dt	<=	119	;
						10'd647	:	dt	<=	130	;
						10'd648	:	dt	<=	139	;
						10'd649	:	dt	<=	145	;
						10'd650	:	dt	<=	171	;
						10'd651	:	dt	<=	174	;
						10'd652	:	dt	<=	182	;
						10'd653	:	dt	<=	159	;
						10'd654	:	dt	<=	193	;
						10'd655	:	dt	<=	150	;
						10'd656	:	dt	<=	137	;
						10'd657	:	dt	<=	110	;
						10'd658	:	dt	<=	84	;
						10'd659	:	dt	<=	78	;
						10'd660	:	dt	<=	75	;
						10'd661	:	dt	<=	162	;
						10'd662	:	dt	<=	190	;
						10'd663	:	dt	<=	191	;
						10'd664	:	dt	<=	193	;
						10'd665	:	dt	<=	193	;
						10'd666	:	dt	<=	194	;
						10'd667	:	dt	<=	195	;
						10'd668	:	dt	<=	195	;
						10'd669	:	dt	<=	195	;
						10'd670	:	dt	<=	194	;
						10'd671	:	dt	<=	194	;
						10'd672	:	dt	<=	92	;
						10'd673	:	dt	<=	107	;
						10'd674	:	dt	<=	120	;
						10'd675	:	dt	<=	130	;
						10'd676	:	dt	<=	138	;
						10'd677	:	dt	<=	146	;
						10'd678	:	dt	<=	162	;
						10'd679	:	dt	<=	192	;
						10'd680	:	dt	<=	174	;
						10'd681	:	dt	<=	154	;
						10'd682	:	dt	<=	180	;
						10'd683	:	dt	<=	137	;
						10'd684	:	dt	<=	117	;
						10'd685	:	dt	<=	95	;
						10'd686	:	dt	<=	79	;
						10'd687	:	dt	<=	75	;
						10'd688	:	dt	<=	82	;
						10'd689	:	dt	<=	176	;
						10'd690	:	dt	<=	191	;
						10'd691	:	dt	<=	192	;
						10'd692	:	dt	<=	193	;
						10'd693	:	dt	<=	194	;
						10'd694	:	dt	<=	195	;
						10'd695	:	dt	<=	195	;
						10'd696	:	dt	<=	196	;
						10'd697	:	dt	<=	196	;
						10'd698	:	dt	<=	195	;
						10'd699	:	dt	<=	195	;
						10'd700	:	dt	<=	90	;
						10'd701	:	dt	<=	107	;
						10'd702	:	dt	<=	120	;
						10'd703	:	dt	<=	129	;
						10'd704	:	dt	<=	137	;
						10'd705	:	dt	<=	146	;
						10'd706	:	dt	<=	156	;
						10'd707	:	dt	<=	186	;
						10'd708	:	dt	<=	167	;
						10'd709	:	dt	<=	146	;
						10'd710	:	dt	<=	159	;
						10'd711	:	dt	<=	127	;
						10'd712	:	dt	<=	105	;
						10'd713	:	dt	<=	90	;
						10'd714	:	dt	<=	79	;
						10'd715	:	dt	<=	71	;
						10'd716	:	dt	<=	96	;
						10'd717	:	dt	<=	184	;
						10'd718	:	dt	<=	190	;
						10'd719	:	dt	<=	193	;
						10'd720	:	dt	<=	194	;
						10'd721	:	dt	<=	195	;
						10'd722	:	dt	<=	196	;
						10'd723	:	dt	<=	196	;
						10'd724	:	dt	<=	196	;
						10'd725	:	dt	<=	196	;
						10'd726	:	dt	<=	195	;
						10'd727	:	dt	<=	195	;
						10'd728	:	dt	<=	89	;
						10'd729	:	dt	<=	106	;
						10'd730	:	dt	<=	117	;
						10'd731	:	dt	<=	127	;
						10'd732	:	dt	<=	136	;
						10'd733	:	dt	<=	145	;
						10'd734	:	dt	<=	151	;
						10'd735	:	dt	<=	171	;
						10'd736	:	dt	<=	156	;
						10'd737	:	dt	<=	148	;
						10'd738	:	dt	<=	151	;
						10'd739	:	dt	<=	133	;
						10'd740	:	dt	<=	117	;
						10'd741	:	dt	<=	98	;
						10'd742	:	dt	<=	80	;
						10'd743	:	dt	<=	68	;
						10'd744	:	dt	<=	108	;
						10'd745	:	dt	<=	186	;
						10'd746	:	dt	<=	189	;
						10'd747	:	dt	<=	190	;
						10'd748	:	dt	<=	193	;
						10'd749	:	dt	<=	193	;
						10'd750	:	dt	<=	194	;
						10'd751	:	dt	<=	194	;
						10'd752	:	dt	<=	195	;
						10'd753	:	dt	<=	195	;
						10'd754	:	dt	<=	195	;
						10'd755	:	dt	<=	195	;
						10'd756	:	dt	<=	89	;
						10'd757	:	dt	<=	106	;
						10'd758	:	dt	<=	116	;
						10'd759	:	dt	<=	127	;
						10'd760	:	dt	<=	136	;
						10'd761	:	dt	<=	145	;
						10'd762	:	dt	<=	151	;
						10'd763	:	dt	<=	163	;
						10'd764	:	dt	<=	159	;
						10'd765	:	dt	<=	154	;
						10'd766	:	dt	<=	152	;
						10'd767	:	dt	<=	144	;
						10'd768	:	dt	<=	129	;
						10'd769	:	dt	<=	100	;
						10'd770	:	dt	<=	78	;
						10'd771	:	dt	<=	64	;
						10'd772	:	dt	<=	115	;
						10'd773	:	dt	<=	186	;
						10'd774	:	dt	<=	187	;
						10'd775	:	dt	<=	189	;
						10'd776	:	dt	<=	192	;
						10'd777	:	dt	<=	193	;
						10'd778	:	dt	<=	194	;
						10'd779	:	dt	<=	194	;
						10'd780	:	dt	<=	194	;
						10'd781	:	dt	<=	195	;
						10'd782	:	dt	<=	195	;
						10'd783	:	dt	<=	194	;
					endcase
				end
				5'd22	:	begin
					case (cnt)
						10'd0	:	dt	<=	186	;
						10'd1	:	dt	<=	187	;
						10'd2	:	dt	<=	188	;
						10'd3	:	dt	<=	186	;
						10'd4	:	dt	<=	188	;
						10'd5	:	dt	<=	189	;
						10'd6	:	dt	<=	188	;
						10'd7	:	dt	<=	188	;
						10'd8	:	dt	<=	187	;
						10'd9	:	dt	<=	189	;
						10'd10	:	dt	<=	189	;
						10'd11	:	dt	<=	188	;
						10'd12	:	dt	<=	187	;
						10'd13	:	dt	<=	185	;
						10'd14	:	dt	<=	184	;
						10'd15	:	dt	<=	181	;
						10'd16	:	dt	<=	183	;
						10'd17	:	dt	<=	183	;
						10'd18	:	dt	<=	181	;
						10'd19	:	dt	<=	178	;
						10'd20	:	dt	<=	177	;
						10'd21	:	dt	<=	176	;
						10'd22	:	dt	<=	174	;
						10'd23	:	dt	<=	172	;
						10'd24	:	dt	<=	169	;
						10'd25	:	dt	<=	167	;
						10'd26	:	dt	<=	164	;
						10'd27	:	dt	<=	161	;
						10'd28	:	dt	<=	191	;
						10'd29	:	dt	<=	191	;
						10'd30	:	dt	<=	191	;
						10'd31	:	dt	<=	191	;
						10'd32	:	dt	<=	192	;
						10'd33	:	dt	<=	193	;
						10'd34	:	dt	<=	193	;
						10'd35	:	dt	<=	191	;
						10'd36	:	dt	<=	191	;
						10'd37	:	dt	<=	192	;
						10'd38	:	dt	<=	198	;
						10'd39	:	dt	<=	194	;
						10'd40	:	dt	<=	190	;
						10'd41	:	dt	<=	189	;
						10'd42	:	dt	<=	191	;
						10'd43	:	dt	<=	192	;
						10'd44	:	dt	<=	186	;
						10'd45	:	dt	<=	186	;
						10'd46	:	dt	<=	183	;
						10'd47	:	dt	<=	182	;
						10'd48	:	dt	<=	182	;
						10'd49	:	dt	<=	181	;
						10'd50	:	dt	<=	177	;
						10'd51	:	dt	<=	175	;
						10'd52	:	dt	<=	173	;
						10'd53	:	dt	<=	171	;
						10'd54	:	dt	<=	169	;
						10'd55	:	dt	<=	166	;
						10'd56	:	dt	<=	195	;
						10'd57	:	dt	<=	195	;
						10'd58	:	dt	<=	195	;
						10'd59	:	dt	<=	196	;
						10'd60	:	dt	<=	197	;
						10'd61	:	dt	<=	196	;
						10'd62	:	dt	<=	196	;
						10'd63	:	dt	<=	195	;
						10'd64	:	dt	<=	195	;
						10'd65	:	dt	<=	198	;
						10'd66	:	dt	<=	160	;
						10'd67	:	dt	<=	188	;
						10'd68	:	dt	<=	197	;
						10'd69	:	dt	<=	194	;
						10'd70	:	dt	<=	180	;
						10'd71	:	dt	<=	168	;
						10'd72	:	dt	<=	192	;
						10'd73	:	dt	<=	189	;
						10'd74	:	dt	<=	187	;
						10'd75	:	dt	<=	187	;
						10'd76	:	dt	<=	184	;
						10'd77	:	dt	<=	183	;
						10'd78	:	dt	<=	181	;
						10'd79	:	dt	<=	178	;
						10'd80	:	dt	<=	179	;
						10'd81	:	dt	<=	178	;
						10'd82	:	dt	<=	171	;
						10'd83	:	dt	<=	170	;
						10'd84	:	dt	<=	197	;
						10'd85	:	dt	<=	198	;
						10'd86	:	dt	<=	200	;
						10'd87	:	dt	<=	200	;
						10'd88	:	dt	<=	200	;
						10'd89	:	dt	<=	200	;
						10'd90	:	dt	<=	201	;
						10'd91	:	dt	<=	200	;
						10'd92	:	dt	<=	198	;
						10'd93	:	dt	<=	196	;
						10'd94	:	dt	<=	129	;
						10'd95	:	dt	<=	146	;
						10'd96	:	dt	<=	207	;
						10'd97	:	dt	<=	197	;
						10'd98	:	dt	<=	194	;
						10'd99	:	dt	<=	110	;
						10'd100	:	dt	<=	179	;
						10'd101	:	dt	<=	196	;
						10'd102	:	dt	<=	191	;
						10'd103	:	dt	<=	191	;
						10'd104	:	dt	<=	190	;
						10'd105	:	dt	<=	187	;
						10'd106	:	dt	<=	183	;
						10'd107	:	dt	<=	186	;
						10'd108	:	dt	<=	148	;
						10'd109	:	dt	<=	160	;
						10'd110	:	dt	<=	179	;
						10'd111	:	dt	<=	172	;
						10'd112	:	dt	<=	201	;
						10'd113	:	dt	<=	201	;
						10'd114	:	dt	<=	203	;
						10'd115	:	dt	<=	203	;
						10'd116	:	dt	<=	202	;
						10'd117	:	dt	<=	203	;
						10'd118	:	dt	<=	203	;
						10'd119	:	dt	<=	203	;
						10'd120	:	dt	<=	201	;
						10'd121	:	dt	<=	194	;
						10'd122	:	dt	<=	154	;
						10'd123	:	dt	<=	109	;
						10'd124	:	dt	<=	207	;
						10'd125	:	dt	<=	198	;
						10'd126	:	dt	<=	204	;
						10'd127	:	dt	<=	110	;
						10'd128	:	dt	<=	152	;
						10'd129	:	dt	<=	205	;
						10'd130	:	dt	<=	193	;
						10'd131	:	dt	<=	193	;
						10'd132	:	dt	<=	192	;
						10'd133	:	dt	<=	189	;
						10'd134	:	dt	<=	187	;
						10'd135	:	dt	<=	196	;
						10'd136	:	dt	<=	119	;
						10'd137	:	dt	<=	111	;
						10'd138	:	dt	<=	189	;
						10'd139	:	dt	<=	173	;
						10'd140	:	dt	<=	204	;
						10'd141	:	dt	<=	204	;
						10'd142	:	dt	<=	207	;
						10'd143	:	dt	<=	208	;
						10'd144	:	dt	<=	205	;
						10'd145	:	dt	<=	206	;
						10'd146	:	dt	<=	208	;
						10'd147	:	dt	<=	206	;
						10'd148	:	dt	<=	204	;
						10'd149	:	dt	<=	203	;
						10'd150	:	dt	<=	177	;
						10'd151	:	dt	<=	91	;
						10'd152	:	dt	<=	192	;
						10'd153	:	dt	<=	204	;
						10'd154	:	dt	<=	205	;
						10'd155	:	dt	<=	110	;
						10'd156	:	dt	<=	127	;
						10'd157	:	dt	<=	211	;
						10'd158	:	dt	<=	195	;
						10'd159	:	dt	<=	196	;
						10'd160	:	dt	<=	193	;
						10'd161	:	dt	<=	190	;
						10'd162	:	dt	<=	195	;
						10'd163	:	dt	<=	190	;
						10'd164	:	dt	<=	98	;
						10'd165	:	dt	<=	123	;
						10'd166	:	dt	<=	192	;
						10'd167	:	dt	<=	179	;
						10'd168	:	dt	<=	206	;
						10'd169	:	dt	<=	208	;
						10'd170	:	dt	<=	210	;
						10'd171	:	dt	<=	211	;
						10'd172	:	dt	<=	209	;
						10'd173	:	dt	<=	209	;
						10'd174	:	dt	<=	211	;
						10'd175	:	dt	<=	209	;
						10'd176	:	dt	<=	210	;
						10'd177	:	dt	<=	203	;
						10'd178	:	dt	<=	180	;
						10'd179	:	dt	<=	85	;
						10'd180	:	dt	<=	170	;
						10'd181	:	dt	<=	214	;
						10'd182	:	dt	<=	207	;
						10'd183	:	dt	<=	118	;
						10'd184	:	dt	<=	115	;
						10'd185	:	dt	<=	211	;
						10'd186	:	dt	<=	198	;
						10'd187	:	dt	<=	199	;
						10'd188	:	dt	<=	198	;
						10'd189	:	dt	<=	193	;
						10'd190	:	dt	<=	202	;
						10'd191	:	dt	<=	170	;
						10'd192	:	dt	<=	84	;
						10'd193	:	dt	<=	150	;
						10'd194	:	dt	<=	193	;
						10'd195	:	dt	<=	181	;
						10'd196	:	dt	<=	211	;
						10'd197	:	dt	<=	212	;
						10'd198	:	dt	<=	211	;
						10'd199	:	dt	<=	212	;
						10'd200	:	dt	<=	212	;
						10'd201	:	dt	<=	212	;
						10'd202	:	dt	<=	213	;
						10'd203	:	dt	<=	212	;
						10'd204	:	dt	<=	213	;
						10'd205	:	dt	<=	209	;
						10'd206	:	dt	<=	193	;
						10'd207	:	dt	<=	114	;
						10'd208	:	dt	<=	137	;
						10'd209	:	dt	<=	222	;
						10'd210	:	dt	<=	213	;
						10'd211	:	dt	<=	132	;
						10'd212	:	dt	<=	104	;
						10'd213	:	dt	<=	210	;
						10'd214	:	dt	<=	202	;
						10'd215	:	dt	<=	204	;
						10'd216	:	dt	<=	199	;
						10'd217	:	dt	<=	198	;
						10'd218	:	dt	<=	208	;
						10'd219	:	dt	<=	145	;
						10'd220	:	dt	<=	83	;
						10'd221	:	dt	<=	182	;
						10'd222	:	dt	<=	188	;
						10'd223	:	dt	<=	184	;
						10'd224	:	dt	<=	214	;
						10'd225	:	dt	<=	213	;
						10'd226	:	dt	<=	213	;
						10'd227	:	dt	<=	215	;
						10'd228	:	dt	<=	215	;
						10'd229	:	dt	<=	216	;
						10'd230	:	dt	<=	215	;
						10'd231	:	dt	<=	213	;
						10'd232	:	dt	<=	214	;
						10'd233	:	dt	<=	214	;
						10'd234	:	dt	<=	207	;
						10'd235	:	dt	<=	144	;
						10'd236	:	dt	<=	108	;
						10'd237	:	dt	<=	221	;
						10'd238	:	dt	<=	215	;
						10'd239	:	dt	<=	121	;
						10'd240	:	dt	<=	90	;
						10'd241	:	dt	<=	209	;
						10'd242	:	dt	<=	205	;
						10'd243	:	dt	<=	205	;
						10'd244	:	dt	<=	200	;
						10'd245	:	dt	<=	207	;
						10'd246	:	dt	<=	200	;
						10'd247	:	dt	<=	124	;
						10'd248	:	dt	<=	104	;
						10'd249	:	dt	<=	202	;
						10'd250	:	dt	<=	189	;
						10'd251	:	dt	<=	187	;
						10'd252	:	dt	<=	217	;
						10'd253	:	dt	<=	216	;
						10'd254	:	dt	<=	216	;
						10'd255	:	dt	<=	217	;
						10'd256	:	dt	<=	218	;
						10'd257	:	dt	<=	217	;
						10'd258	:	dt	<=	218	;
						10'd259	:	dt	<=	217	;
						10'd260	:	dt	<=	218	;
						10'd261	:	dt	<=	218	;
						10'd262	:	dt	<=	213	;
						10'd263	:	dt	<=	158	;
						10'd264	:	dt	<=	79	;
						10'd265	:	dt	<=	209	;
						10'd266	:	dt	<=	219	;
						10'd267	:	dt	<=	116	;
						10'd268	:	dt	<=	88	;
						10'd269	:	dt	<=	206	;
						10'd270	:	dt	<=	210	;
						10'd271	:	dt	<=	207	;
						10'd272	:	dt	<=	203	;
						10'd273	:	dt	<=	205	;
						10'd274	:	dt	<=	175	;
						10'd275	:	dt	<=	88	;
						10'd276	:	dt	<=	146	;
						10'd277	:	dt	<=	205	;
						10'd278	:	dt	<=	191	;
						10'd279	:	dt	<=	191	;
						10'd280	:	dt	<=	218	;
						10'd281	:	dt	<=	219	;
						10'd282	:	dt	<=	219	;
						10'd283	:	dt	<=	219	;
						10'd284	:	dt	<=	220	;
						10'd285	:	dt	<=	219	;
						10'd286	:	dt	<=	218	;
						10'd287	:	dt	<=	219	;
						10'd288	:	dt	<=	220	;
						10'd289	:	dt	<=	220	;
						10'd290	:	dt	<=	212	;
						10'd291	:	dt	<=	180	;
						10'd292	:	dt	<=	84	;
						10'd293	:	dt	<=	167	;
						10'd294	:	dt	<=	228	;
						10'd295	:	dt	<=	133	;
						10'd296	:	dt	<=	92	;
						10'd297	:	dt	<=	203	;
						10'd298	:	dt	<=	215	;
						10'd299	:	dt	<=	208	;
						10'd300	:	dt	<=	206	;
						10'd301	:	dt	<=	194	;
						10'd302	:	dt	<=	141	;
						10'd303	:	dt	<=	73	;
						10'd304	:	dt	<=	193	;
						10'd305	:	dt	<=	199	;
						10'd306	:	dt	<=	193	;
						10'd307	:	dt	<=	192	;
						10'd308	:	dt	<=	220	;
						10'd309	:	dt	<=	220	;
						10'd310	:	dt	<=	220	;
						10'd311	:	dt	<=	220	;
						10'd312	:	dt	<=	221	;
						10'd313	:	dt	<=	220	;
						10'd314	:	dt	<=	220	;
						10'd315	:	dt	<=	221	;
						10'd316	:	dt	<=	220	;
						10'd317	:	dt	<=	223	;
						10'd318	:	dt	<=	205	;
						10'd319	:	dt	<=	188	;
						10'd320	:	dt	<=	137	;
						10'd321	:	dt	<=	104	;
						10'd322	:	dt	<=	218	;
						10'd323	:	dt	<=	141	;
						10'd324	:	dt	<=	88	;
						10'd325	:	dt	<=	201	;
						10'd326	:	dt	<=	220	;
						10'd327	:	dt	<=	211	;
						10'd328	:	dt	<=	213	;
						10'd329	:	dt	<=	200	;
						10'd330	:	dt	<=	112	;
						10'd331	:	dt	<=	114	;
						10'd332	:	dt	<=	215	;
						10'd333	:	dt	<=	197	;
						10'd334	:	dt	<=	198	;
						10'd335	:	dt	<=	195	;
						10'd336	:	dt	<=	223	;
						10'd337	:	dt	<=	222	;
						10'd338	:	dt	<=	222	;
						10'd339	:	dt	<=	222	;
						10'd340	:	dt	<=	222	;
						10'd341	:	dt	<=	222	;
						10'd342	:	dt	<=	222	;
						10'd343	:	dt	<=	223	;
						10'd344	:	dt	<=	222	;
						10'd345	:	dt	<=	224	;
						10'd346	:	dt	<=	215	;
						10'd347	:	dt	<=	195	;
						10'd348	:	dt	<=	169	;
						10'd349	:	dt	<=	123	;
						10'd350	:	dt	<=	180	;
						10'd351	:	dt	<=	143	;
						10'd352	:	dt	<=	108	;
						10'd353	:	dt	<=	169	;
						10'd354	:	dt	<=	222	;
						10'd355	:	dt	<=	216	;
						10'd356	:	dt	<=	208	;
						10'd357	:	dt	<=	178	;
						10'd358	:	dt	<=	88	;
						10'd359	:	dt	<=	172	;
						10'd360	:	dt	<=	214	;
						10'd361	:	dt	<=	201	;
						10'd362	:	dt	<=	201	;
						10'd363	:	dt	<=	200	;
						10'd364	:	dt	<=	225	;
						10'd365	:	dt	<=	225	;
						10'd366	:	dt	<=	225	;
						10'd367	:	dt	<=	225	;
						10'd368	:	dt	<=	224	;
						10'd369	:	dt	<=	225	;
						10'd370	:	dt	<=	225	;
						10'd371	:	dt	<=	225	;
						10'd372	:	dt	<=	224	;
						10'd373	:	dt	<=	226	;
						10'd374	:	dt	<=	226	;
						10'd375	:	dt	<=	200	;
						10'd376	:	dt	<=	197	;
						10'd377	:	dt	<=	211	;
						10'd378	:	dt	<=	203	;
						10'd379	:	dt	<=	180	;
						10'd380	:	dt	<=	188	;
						10'd381	:	dt	<=	113	;
						10'd382	:	dt	<=	118	;
						10'd383	:	dt	<=	199	;
						10'd384	:	dt	<=	199	;
						10'd385	:	dt	<=	135	;
						10'd386	:	dt	<=	91	;
						10'd387	:	dt	<=	211	;
						10'd388	:	dt	<=	207	;
						10'd389	:	dt	<=	203	;
						10'd390	:	dt	<=	202	;
						10'd391	:	dt	<=	199	;
						10'd392	:	dt	<=	227	;
						10'd393	:	dt	<=	227	;
						10'd394	:	dt	<=	227	;
						10'd395	:	dt	<=	227	;
						10'd396	:	dt	<=	227	;
						10'd397	:	dt	<=	227	;
						10'd398	:	dt	<=	226	;
						10'd399	:	dt	<=	226	;
						10'd400	:	dt	<=	227	;
						10'd401	:	dt	<=	227	;
						10'd402	:	dt	<=	230	;
						10'd403	:	dt	<=	213	;
						10'd404	:	dt	<=	201	;
						10'd405	:	dt	<=	181	;
						10'd406	:	dt	<=	168	;
						10'd407	:	dt	<=	172	;
						10'd408	:	dt	<=	185	;
						10'd409	:	dt	<=	120	;
						10'd410	:	dt	<=	72	;
						10'd411	:	dt	<=	84	;
						10'd412	:	dt	<=	128	;
						10'd413	:	dt	<=	83	;
						10'd414	:	dt	<=	138	;
						10'd415	:	dt	<=	225	;
						10'd416	:	dt	<=	206	;
						10'd417	:	dt	<=	205	;
						10'd418	:	dt	<=	204	;
						10'd419	:	dt	<=	200	;
						10'd420	:	dt	<=	228	;
						10'd421	:	dt	<=	228	;
						10'd422	:	dt	<=	228	;
						10'd423	:	dt	<=	228	;
						10'd424	:	dt	<=	227	;
						10'd425	:	dt	<=	228	;
						10'd426	:	dt	<=	229	;
						10'd427	:	dt	<=	229	;
						10'd428	:	dt	<=	230	;
						10'd429	:	dt	<=	228	;
						10'd430	:	dt	<=	229	;
						10'd431	:	dt	<=	224	;
						10'd432	:	dt	<=	214	;
						10'd433	:	dt	<=	150	;
						10'd434	:	dt	<=	56	;
						10'd435	:	dt	<=	99	;
						10'd436	:	dt	<=	175	;
						10'd437	:	dt	<=	142	;
						10'd438	:	dt	<=	108	;
						10'd439	:	dt	<=	94	;
						10'd440	:	dt	<=	95	;
						10'd441	:	dt	<=	49	;
						10'd442	:	dt	<=	183	;
						10'd443	:	dt	<=	221	;
						10'd444	:	dt	<=	211	;
						10'd445	:	dt	<=	209	;
						10'd446	:	dt	<=	206	;
						10'd447	:	dt	<=	203	;
						10'd448	:	dt	<=	229	;
						10'd449	:	dt	<=	230	;
						10'd450	:	dt	<=	230	;
						10'd451	:	dt	<=	230	;
						10'd452	:	dt	<=	229	;
						10'd453	:	dt	<=	229	;
						10'd454	:	dt	<=	230	;
						10'd455	:	dt	<=	230	;
						10'd456	:	dt	<=	230	;
						10'd457	:	dt	<=	230	;
						10'd458	:	dt	<=	229	;
						10'd459	:	dt	<=	225	;
						10'd460	:	dt	<=	201	;
						10'd461	:	dt	<=	125	;
						10'd462	:	dt	<=	70	;
						10'd463	:	dt	<=	41	;
						10'd464	:	dt	<=	118	;
						10'd465	:	dt	<=	151	;
						10'd466	:	dt	<=	128	;
						10'd467	:	dt	<=	120	;
						10'd468	:	dt	<=	116	;
						10'd469	:	dt	<=	42	;
						10'd470	:	dt	<=	191	;
						10'd471	:	dt	<=	223	;
						10'd472	:	dt	<=	213	;
						10'd473	:	dt	<=	212	;
						10'd474	:	dt	<=	209	;
						10'd475	:	dt	<=	206	;
						10'd476	:	dt	<=	231	;
						10'd477	:	dt	<=	231	;
						10'd478	:	dt	<=	231	;
						10'd479	:	dt	<=	231	;
						10'd480	:	dt	<=	232	;
						10'd481	:	dt	<=	231	;
						10'd482	:	dt	<=	231	;
						10'd483	:	dt	<=	232	;
						10'd484	:	dt	<=	232	;
						10'd485	:	dt	<=	231	;
						10'd486	:	dt	<=	231	;
						10'd487	:	dt	<=	221	;
						10'd488	:	dt	<=	198	;
						10'd489	:	dt	<=	161	;
						10'd490	:	dt	<=	110	;
						10'd491	:	dt	<=	55	;
						10'd492	:	dt	<=	50	;
						10'd493	:	dt	<=	61	;
						10'd494	:	dt	<=	98	;
						10'd495	:	dt	<=	121	;
						10'd496	:	dt	<=	91	;
						10'd497	:	dt	<=	35	;
						10'd498	:	dt	<=	142	;
						10'd499	:	dt	<=	233	;
						10'd500	:	dt	<=	212	;
						10'd501	:	dt	<=	214	;
						10'd502	:	dt	<=	209	;
						10'd503	:	dt	<=	208	;
						10'd504	:	dt	<=	234	;
						10'd505	:	dt	<=	233	;
						10'd506	:	dt	<=	235	;
						10'd507	:	dt	<=	234	;
						10'd508	:	dt	<=	235	;
						10'd509	:	dt	<=	235	;
						10'd510	:	dt	<=	235	;
						10'd511	:	dt	<=	235	;
						10'd512	:	dt	<=	236	;
						10'd513	:	dt	<=	235	;
						10'd514	:	dt	<=	233	;
						10'd515	:	dt	<=	215	;
						10'd516	:	dt	<=	203	;
						10'd517	:	dt	<=	171	;
						10'd518	:	dt	<=	102	;
						10'd519	:	dt	<=	59	;
						10'd520	:	dt	<=	67	;
						10'd521	:	dt	<=	69	;
						10'd522	:	dt	<=	102	;
						10'd523	:	dt	<=	163	;
						10'd524	:	dt	<=	126	;
						10'd525	:	dt	<=	65	;
						10'd526	:	dt	<=	73	;
						10'd527	:	dt	<=	226	;
						10'd528	:	dt	<=	214	;
						10'd529	:	dt	<=	214	;
						10'd530	:	dt	<=	211	;
						10'd531	:	dt	<=	210	;
						10'd532	:	dt	<=	235	;
						10'd533	:	dt	<=	235	;
						10'd534	:	dt	<=	236	;
						10'd535	:	dt	<=	236	;
						10'd536	:	dt	<=	236	;
						10'd537	:	dt	<=	237	;
						10'd538	:	dt	<=	236	;
						10'd539	:	dt	<=	237	;
						10'd540	:	dt	<=	238	;
						10'd541	:	dt	<=	238	;
						10'd542	:	dt	<=	234	;
						10'd543	:	dt	<=	213	;
						10'd544	:	dt	<=	203	;
						10'd545	:	dt	<=	156	;
						10'd546	:	dt	<=	103	;
						10'd547	:	dt	<=	73	;
						10'd548	:	dt	<=	75	;
						10'd549	:	dt	<=	111	;
						10'd550	:	dt	<=	190	;
						10'd551	:	dt	<=	201	;
						10'd552	:	dt	<=	169	;
						10'd553	:	dt	<=	111	;
						10'd554	:	dt	<=	35	;
						10'd555	:	dt	<=	158	;
						10'd556	:	dt	<=	229	;
						10'd557	:	dt	<=	213	;
						10'd558	:	dt	<=	213	;
						10'd559	:	dt	<=	211	;
						10'd560	:	dt	<=	235	;
						10'd561	:	dt	<=	234	;
						10'd562	:	dt	<=	235	;
						10'd563	:	dt	<=	236	;
						10'd564	:	dt	<=	236	;
						10'd565	:	dt	<=	236	;
						10'd566	:	dt	<=	237	;
						10'd567	:	dt	<=	237	;
						10'd568	:	dt	<=	238	;
						10'd569	:	dt	<=	237	;
						10'd570	:	dt	<=	235	;
						10'd571	:	dt	<=	216	;
						10'd572	:	dt	<=	205	;
						10'd573	:	dt	<=	175	;
						10'd574	:	dt	<=	124	;
						10'd575	:	dt	<=	80	;
						10'd576	:	dt	<=	82	;
						10'd577	:	dt	<=	152	;
						10'd578	:	dt	<=	217	;
						10'd579	:	dt	<=	226	;
						10'd580	:	dt	<=	196	;
						10'd581	:	dt	<=	155	;
						10'd582	:	dt	<=	48	;
						10'd583	:	dt	<=	111	;
						10'd584	:	dt	<=	235	;
						10'd585	:	dt	<=	212	;
						10'd586	:	dt	<=	214	;
						10'd587	:	dt	<=	211	;
						10'd588	:	dt	<=	235	;
						10'd589	:	dt	<=	234	;
						10'd590	:	dt	<=	236	;
						10'd591	:	dt	<=	236	;
						10'd592	:	dt	<=	235	;
						10'd593	:	dt	<=	236	;
						10'd594	:	dt	<=	237	;
						10'd595	:	dt	<=	237	;
						10'd596	:	dt	<=	237	;
						10'd597	:	dt	<=	236	;
						10'd598	:	dt	<=	236	;
						10'd599	:	dt	<=	213	;
						10'd600	:	dt	<=	203	;
						10'd601	:	dt	<=	183	;
						10'd602	:	dt	<=	134	;
						10'd603	:	dt	<=	80	;
						10'd604	:	dt	<=	94	;
						10'd605	:	dt	<=	178	;
						10'd606	:	dt	<=	223	;
						10'd607	:	dt	<=	218	;
						10'd608	:	dt	<=	191	;
						10'd609	:	dt	<=	138	;
						10'd610	:	dt	<=	41	;
						10'd611	:	dt	<=	131	;
						10'd612	:	dt	<=	232	;
						10'd613	:	dt	<=	210	;
						10'd614	:	dt	<=	212	;
						10'd615	:	dt	<=	211	;
						10'd616	:	dt	<=	236	;
						10'd617	:	dt	<=	236	;
						10'd618	:	dt	<=	237	;
						10'd619	:	dt	<=	237	;
						10'd620	:	dt	<=	237	;
						10'd621	:	dt	<=	238	;
						10'd622	:	dt	<=	238	;
						10'd623	:	dt	<=	238	;
						10'd624	:	dt	<=	239	;
						10'd625	:	dt	<=	238	;
						10'd626	:	dt	<=	238	;
						10'd627	:	dt	<=	208	;
						10'd628	:	dt	<=	195	;
						10'd629	:	dt	<=	200	;
						10'd630	:	dt	<=	140	;
						10'd631	:	dt	<=	88	;
						10'd632	:	dt	<=	106	;
						10'd633	:	dt	<=	199	;
						10'd634	:	dt	<=	227	;
						10'd635	:	dt	<=	198	;
						10'd636	:	dt	<=	158	;
						10'd637	:	dt	<=	111	;
						10'd638	:	dt	<=	29	;
						10'd639	:	dt	<=	173	;
						10'd640	:	dt	<=	225	;
						10'd641	:	dt	<=	211	;
						10'd642	:	dt	<=	212	;
						10'd643	:	dt	<=	208	;
						10'd644	:	dt	<=	238	;
						10'd645	:	dt	<=	238	;
						10'd646	:	dt	<=	238	;
						10'd647	:	dt	<=	238	;
						10'd648	:	dt	<=	239	;
						10'd649	:	dt	<=	239	;
						10'd650	:	dt	<=	239	;
						10'd651	:	dt	<=	240	;
						10'd652	:	dt	<=	240	;
						10'd653	:	dt	<=	239	;
						10'd654	:	dt	<=	239	;
						10'd655	:	dt	<=	203	;
						10'd656	:	dt	<=	190	;
						10'd657	:	dt	<=	194	;
						10'd658	:	dt	<=	143	;
						10'd659	:	dt	<=	92	;
						10'd660	:	dt	<=	105	;
						10'd661	:	dt	<=	211	;
						10'd662	:	dt	<=	210	;
						10'd663	:	dt	<=	175	;
						10'd664	:	dt	<=	130	;
						10'd665	:	dt	<=	94	;
						10'd666	:	dt	<=	47	;
						10'd667	:	dt	<=	207	;
						10'd668	:	dt	<=	221	;
						10'd669	:	dt	<=	214	;
						10'd670	:	dt	<=	215	;
						10'd671	:	dt	<=	220	;
						10'd672	:	dt	<=	237	;
						10'd673	:	dt	<=	238	;
						10'd674	:	dt	<=	238	;
						10'd675	:	dt	<=	237	;
						10'd676	:	dt	<=	237	;
						10'd677	:	dt	<=	238	;
						10'd678	:	dt	<=	239	;
						10'd679	:	dt	<=	239	;
						10'd680	:	dt	<=	239	;
						10'd681	:	dt	<=	239	;
						10'd682	:	dt	<=	241	;
						10'd683	:	dt	<=	202	;
						10'd684	:	dt	<=	183	;
						10'd685	:	dt	<=	181	;
						10'd686	:	dt	<=	144	;
						10'd687	:	dt	<=	89	;
						10'd688	:	dt	<=	92	;
						10'd689	:	dt	<=	192	;
						10'd690	:	dt	<=	190	;
						10'd691	:	dt	<=	170	;
						10'd692	:	dt	<=	119	;
						10'd693	:	dt	<=	70	;
						10'd694	:	dt	<=	68	;
						10'd695	:	dt	<=	222	;
						10'd696	:	dt	<=	219	;
						10'd697	:	dt	<=	227	;
						10'd698	:	dt	<=	214	;
						10'd699	:	dt	<=	145	;
						10'd700	:	dt	<=	244	;
						10'd701	:	dt	<=	247	;
						10'd702	:	dt	<=	248	;
						10'd703	:	dt	<=	248	;
						10'd704	:	dt	<=	248	;
						10'd705	:	dt	<=	249	;
						10'd706	:	dt	<=	251	;
						10'd707	:	dt	<=	250	;
						10'd708	:	dt	<=	250	;
						10'd709	:	dt	<=	247	;
						10'd710	:	dt	<=	252	;
						10'd711	:	dt	<=	220	;
						10'd712	:	dt	<=	181	;
						10'd713	:	dt	<=	182	;
						10'd714	:	dt	<=	143	;
						10'd715	:	dt	<=	97	;
						10'd716	:	dt	<=	94	;
						10'd717	:	dt	<=	184	;
						10'd718	:	dt	<=	186	;
						10'd719	:	dt	<=	155	;
						10'd720	:	dt	<=	100	;
						10'd721	:	dt	<=	38	;
						10'd722	:	dt	<=	113	;
						10'd723	:	dt	<=	247	;
						10'd724	:	dt	<=	214	;
						10'd725	:	dt	<=	157	;
						10'd726	:	dt	<=	82	;
						10'd727	:	dt	<=	24	;
						10'd728	:	dt	<=	151	;
						10'd729	:	dt	<=	156	;
						10'd730	:	dt	<=	161	;
						10'd731	:	dt	<=	169	;
						10'd732	:	dt	<=	174	;
						10'd733	:	dt	<=	178	;
						10'd734	:	dt	<=	184	;
						10'd735	:	dt	<=	186	;
						10'd736	:	dt	<=	191	;
						10'd737	:	dt	<=	198	;
						10'd738	:	dt	<=	205	;
						10'd739	:	dt	<=	202	;
						10'd740	:	dt	<=	182	;
						10'd741	:	dt	<=	173	;
						10'd742	:	dt	<=	141	;
						10'd743	:	dt	<=	117	;
						10'd744	:	dt	<=	90	;
						10'd745	:	dt	<=	170	;
						10'd746	:	dt	<=	177	;
						10'd747	:	dt	<=	130	;
						10'd748	:	dt	<=	76	;
						10'd749	:	dt	<=	30	;
						10'd750	:	dt	<=	150	;
						10'd751	:	dt	<=	159	;
						10'd752	:	dt	<=	73	;
						10'd753	:	dt	<=	27	;
						10'd754	:	dt	<=	24	;
						10'd755	:	dt	<=	21	;
						10'd756	:	dt	<=	94	;
						10'd757	:	dt	<=	93	;
						10'd758	:	dt	<=	94	;
						10'd759	:	dt	<=	96	;
						10'd760	:	dt	<=	94	;
						10'd761	:	dt	<=	93	;
						10'd762	:	dt	<=	94	;
						10'd763	:	dt	<=	92	;
						10'd764	:	dt	<=	91	;
						10'd765	:	dt	<=	95	;
						10'd766	:	dt	<=	93	;
						10'd767	:	dt	<=	109	;
						10'd768	:	dt	<=	189	;
						10'd769	:	dt	<=	174	;
						10'd770	:	dt	<=	140	;
						10'd771	:	dt	<=	120	;
						10'd772	:	dt	<=	82	;
						10'd773	:	dt	<=	127	;
						10'd774	:	dt	<=	135	;
						10'd775	:	dt	<=	85	;
						10'd776	:	dt	<=	47	;
						10'd777	:	dt	<=	28	;
						10'd778	:	dt	<=	48	;
						10'd779	:	dt	<=	31	;
						10'd780	:	dt	<=	6	;
						10'd781	:	dt	<=	19	;
						10'd782	:	dt	<=	32	;
						10'd783	:	dt	<=	13	;
					endcase
				end
				5'd23	:	begin
					case (cnt)
						10'd0	:	dt	<=	119	;
						10'd1	:	dt	<=	122	;
						10'd2	:	dt	<=	125	;
						10'd3	:	dt	<=	134	;
						10'd4	:	dt	<=	144	;
						10'd5	:	dt	<=	154	;
						10'd6	:	dt	<=	161	;
						10'd7	:	dt	<=	164	;
						10'd8	:	dt	<=	167	;
						10'd9	:	dt	<=	171	;
						10'd10	:	dt	<=	177	;
						10'd11	:	dt	<=	181	;
						10'd12	:	dt	<=	184	;
						10'd13	:	dt	<=	187	;
						10'd14	:	dt	<=	189	;
						10'd15	:	dt	<=	191	;
						10'd16	:	dt	<=	194	;
						10'd17	:	dt	<=	196	;
						10'd18	:	dt	<=	198	;
						10'd19	:	dt	<=	198	;
						10'd20	:	dt	<=	197	;
						10'd21	:	dt	<=	198	;
						10'd22	:	dt	<=	198	;
						10'd23	:	dt	<=	199	;
						10'd24	:	dt	<=	200	;
						10'd25	:	dt	<=	199	;
						10'd26	:	dt	<=	198	;
						10'd27	:	dt	<=	198	;
						10'd28	:	dt	<=	119	;
						10'd29	:	dt	<=	122	;
						10'd30	:	dt	<=	127	;
						10'd31	:	dt	<=	136	;
						10'd32	:	dt	<=	146	;
						10'd33	:	dt	<=	155	;
						10'd34	:	dt	<=	162	;
						10'd35	:	dt	<=	166	;
						10'd36	:	dt	<=	168	;
						10'd37	:	dt	<=	174	;
						10'd38	:	dt	<=	179	;
						10'd39	:	dt	<=	183	;
						10'd40	:	dt	<=	187	;
						10'd41	:	dt	<=	188	;
						10'd42	:	dt	<=	189	;
						10'd43	:	dt	<=	192	;
						10'd44	:	dt	<=	197	;
						10'd45	:	dt	<=	198	;
						10'd46	:	dt	<=	198	;
						10'd47	:	dt	<=	200	;
						10'd48	:	dt	<=	200	;
						10'd49	:	dt	<=	200	;
						10'd50	:	dt	<=	200	;
						10'd51	:	dt	<=	201	;
						10'd52	:	dt	<=	201	;
						10'd53	:	dt	<=	200	;
						10'd54	:	dt	<=	199	;
						10'd55	:	dt	<=	199	;
						10'd56	:	dt	<=	120	;
						10'd57	:	dt	<=	123	;
						10'd58	:	dt	<=	127	;
						10'd59	:	dt	<=	137	;
						10'd60	:	dt	<=	147	;
						10'd61	:	dt	<=	157	;
						10'd62	:	dt	<=	164	;
						10'd63	:	dt	<=	167	;
						10'd64	:	dt	<=	169	;
						10'd65	:	dt	<=	175	;
						10'd66	:	dt	<=	180	;
						10'd67	:	dt	<=	184	;
						10'd68	:	dt	<=	188	;
						10'd69	:	dt	<=	190	;
						10'd70	:	dt	<=	192	;
						10'd71	:	dt	<=	195	;
						10'd72	:	dt	<=	197	;
						10'd73	:	dt	<=	199	;
						10'd74	:	dt	<=	201	;
						10'd75	:	dt	<=	202	;
						10'd76	:	dt	<=	202	;
						10'd77	:	dt	<=	203	;
						10'd78	:	dt	<=	203	;
						10'd79	:	dt	<=	202	;
						10'd80	:	dt	<=	202	;
						10'd81	:	dt	<=	202	;
						10'd82	:	dt	<=	201	;
						10'd83	:	dt	<=	201	;
						10'd84	:	dt	<=	120	;
						10'd85	:	dt	<=	123	;
						10'd86	:	dt	<=	127	;
						10'd87	:	dt	<=	138	;
						10'd88	:	dt	<=	148	;
						10'd89	:	dt	<=	158	;
						10'd90	:	dt	<=	165	;
						10'd91	:	dt	<=	168	;
						10'd92	:	dt	<=	170	;
						10'd93	:	dt	<=	176	;
						10'd94	:	dt	<=	182	;
						10'd95	:	dt	<=	186	;
						10'd96	:	dt	<=	189	;
						10'd97	:	dt	<=	192	;
						10'd98	:	dt	<=	195	;
						10'd99	:	dt	<=	196	;
						10'd100	:	dt	<=	198	;
						10'd101	:	dt	<=	201	;
						10'd102	:	dt	<=	203	;
						10'd103	:	dt	<=	203	;
						10'd104	:	dt	<=	203	;
						10'd105	:	dt	<=	203	;
						10'd106	:	dt	<=	203	;
						10'd107	:	dt	<=	203	;
						10'd108	:	dt	<=	203	;
						10'd109	:	dt	<=	203	;
						10'd110	:	dt	<=	203	;
						10'd111	:	dt	<=	202	;
						10'd112	:	dt	<=	122	;
						10'd113	:	dt	<=	124	;
						10'd114	:	dt	<=	127	;
						10'd115	:	dt	<=	138	;
						10'd116	:	dt	<=	149	;
						10'd117	:	dt	<=	159	;
						10'd118	:	dt	<=	166	;
						10'd119	:	dt	<=	169	;
						10'd120	:	dt	<=	173	;
						10'd121	:	dt	<=	178	;
						10'd122	:	dt	<=	183	;
						10'd123	:	dt	<=	188	;
						10'd124	:	dt	<=	190	;
						10'd125	:	dt	<=	192	;
						10'd126	:	dt	<=	196	;
						10'd127	:	dt	<=	197	;
						10'd128	:	dt	<=	200	;
						10'd129	:	dt	<=	202	;
						10'd130	:	dt	<=	202	;
						10'd131	:	dt	<=	203	;
						10'd132	:	dt	<=	204	;
						10'd133	:	dt	<=	203	;
						10'd134	:	dt	<=	204	;
						10'd135	:	dt	<=	203	;
						10'd136	:	dt	<=	204	;
						10'd137	:	dt	<=	204	;
						10'd138	:	dt	<=	204	;
						10'd139	:	dt	<=	201	;
						10'd140	:	dt	<=	121	;
						10'd141	:	dt	<=	124	;
						10'd142	:	dt	<=	129	;
						10'd143	:	dt	<=	140	;
						10'd144	:	dt	<=	150	;
						10'd145	:	dt	<=	160	;
						10'd146	:	dt	<=	166	;
						10'd147	:	dt	<=	170	;
						10'd148	:	dt	<=	174	;
						10'd149	:	dt	<=	179	;
						10'd150	:	dt	<=	184	;
						10'd151	:	dt	<=	189	;
						10'd152	:	dt	<=	191	;
						10'd153	:	dt	<=	194	;
						10'd154	:	dt	<=	197	;
						10'd155	:	dt	<=	199	;
						10'd156	:	dt	<=	201	;
						10'd157	:	dt	<=	203	;
						10'd158	:	dt	<=	203	;
						10'd159	:	dt	<=	204	;
						10'd160	:	dt	<=	207	;
						10'd161	:	dt	<=	206	;
						10'd162	:	dt	<=	205	;
						10'd163	:	dt	<=	205	;
						10'd164	:	dt	<=	204	;
						10'd165	:	dt	<=	204	;
						10'd166	:	dt	<=	204	;
						10'd167	:	dt	<=	203	;
						10'd168	:	dt	<=	121	;
						10'd169	:	dt	<=	123	;
						10'd170	:	dt	<=	129	;
						10'd171	:	dt	<=	141	;
						10'd172	:	dt	<=	151	;
						10'd173	:	dt	<=	161	;
						10'd174	:	dt	<=	168	;
						10'd175	:	dt	<=	169	;
						10'd176	:	dt	<=	174	;
						10'd177	:	dt	<=	180	;
						10'd178	:	dt	<=	186	;
						10'd179	:	dt	<=	190	;
						10'd180	:	dt	<=	193	;
						10'd181	:	dt	<=	196	;
						10'd182	:	dt	<=	199	;
						10'd183	:	dt	<=	201	;
						10'd184	:	dt	<=	203	;
						10'd185	:	dt	<=	203	;
						10'd186	:	dt	<=	206	;
						10'd187	:	dt	<=	206	;
						10'd188	:	dt	<=	204	;
						10'd189	:	dt	<=	205	;
						10'd190	:	dt	<=	203	;
						10'd191	:	dt	<=	206	;
						10'd192	:	dt	<=	208	;
						10'd193	:	dt	<=	205	;
						10'd194	:	dt	<=	203	;
						10'd195	:	dt	<=	204	;
						10'd196	:	dt	<=	122	;
						10'd197	:	dt	<=	124	;
						10'd198	:	dt	<=	130	;
						10'd199	:	dt	<=	142	;
						10'd200	:	dt	<=	152	;
						10'd201	:	dt	<=	162	;
						10'd202	:	dt	<=	169	;
						10'd203	:	dt	<=	172	;
						10'd204	:	dt	<=	175	;
						10'd205	:	dt	<=	182	;
						10'd206	:	dt	<=	187	;
						10'd207	:	dt	<=	191	;
						10'd208	:	dt	<=	195	;
						10'd209	:	dt	<=	197	;
						10'd210	:	dt	<=	200	;
						10'd211	:	dt	<=	203	;
						10'd212	:	dt	<=	203	;
						10'd213	:	dt	<=	206	;
						10'd214	:	dt	<=	206	;
						10'd215	:	dt	<=	203	;
						10'd216	:	dt	<=	230	;
						10'd217	:	dt	<=	238	;
						10'd218	:	dt	<=	214	;
						10'd219	:	dt	<=	207	;
						10'd220	:	dt	<=	203	;
						10'd221	:	dt	<=	205	;
						10'd222	:	dt	<=	206	;
						10'd223	:	dt	<=	204	;
						10'd224	:	dt	<=	121	;
						10'd225	:	dt	<=	124	;
						10'd226	:	dt	<=	131	;
						10'd227	:	dt	<=	143	;
						10'd228	:	dt	<=	152	;
						10'd229	:	dt	<=	162	;
						10'd230	:	dt	<=	169	;
						10'd231	:	dt	<=	172	;
						10'd232	:	dt	<=	176	;
						10'd233	:	dt	<=	183	;
						10'd234	:	dt	<=	189	;
						10'd235	:	dt	<=	193	;
						10'd236	:	dt	<=	196	;
						10'd237	:	dt	<=	198	;
						10'd238	:	dt	<=	202	;
						10'd239	:	dt	<=	204	;
						10'd240	:	dt	<=	206	;
						10'd241	:	dt	<=	206	;
						10'd242	:	dt	<=	210	;
						10'd243	:	dt	<=	247	;
						10'd244	:	dt	<=	255	;
						10'd245	:	dt	<=	224	;
						10'd246	:	dt	<=	220	;
						10'd247	:	dt	<=	197	;
						10'd248	:	dt	<=	142	;
						10'd249	:	dt	<=	200	;
						10'd250	:	dt	<=	210	;
						10'd251	:	dt	<=	207	;
						10'd252	:	dt	<=	122	;
						10'd253	:	dt	<=	124	;
						10'd254	:	dt	<=	131	;
						10'd255	:	dt	<=	143	;
						10'd256	:	dt	<=	154	;
						10'd257	:	dt	<=	164	;
						10'd258	:	dt	<=	171	;
						10'd259	:	dt	<=	174	;
						10'd260	:	dt	<=	178	;
						10'd261	:	dt	<=	185	;
						10'd262	:	dt	<=	191	;
						10'd263	:	dt	<=	194	;
						10'd264	:	dt	<=	197	;
						10'd265	:	dt	<=	201	;
						10'd266	:	dt	<=	203	;
						10'd267	:	dt	<=	206	;
						10'd268	:	dt	<=	205	;
						10'd269	:	dt	<=	215	;
						10'd270	:	dt	<=	255	;
						10'd271	:	dt	<=	240	;
						10'd272	:	dt	<=	204	;
						10'd273	:	dt	<=	143	;
						10'd274	:	dt	<=	171	;
						10'd275	:	dt	<=	178	;
						10'd276	:	dt	<=	181	;
						10'd277	:	dt	<=	211	;
						10'd278	:	dt	<=	209	;
						10'd279	:	dt	<=	209	;
						10'd280	:	dt	<=	122	;
						10'd281	:	dt	<=	125	;
						10'd282	:	dt	<=	132	;
						10'd283	:	dt	<=	144	;
						10'd284	:	dt	<=	155	;
						10'd285	:	dt	<=	165	;
						10'd286	:	dt	<=	172	;
						10'd287	:	dt	<=	174	;
						10'd288	:	dt	<=	179	;
						10'd289	:	dt	<=	186	;
						10'd290	:	dt	<=	191	;
						10'd291	:	dt	<=	196	;
						10'd292	:	dt	<=	199	;
						10'd293	:	dt	<=	201	;
						10'd294	:	dt	<=	203	;
						10'd295	:	dt	<=	208	;
						10'd296	:	dt	<=	203	;
						10'd297	:	dt	<=	249	;
						10'd298	:	dt	<=	255	;
						10'd299	:	dt	<=	167	;
						10'd300	:	dt	<=	122	;
						10'd301	:	dt	<=	184	;
						10'd302	:	dt	<=	213	;
						10'd303	:	dt	<=	213	;
						10'd304	:	dt	<=	217	;
						10'd305	:	dt	<=	212	;
						10'd306	:	dt	<=	210	;
						10'd307	:	dt	<=	210	;
						10'd308	:	dt	<=	122	;
						10'd309	:	dt	<=	124	;
						10'd310	:	dt	<=	132	;
						10'd311	:	dt	<=	145	;
						10'd312	:	dt	<=	156	;
						10'd313	:	dt	<=	167	;
						10'd314	:	dt	<=	173	;
						10'd315	:	dt	<=	175	;
						10'd316	:	dt	<=	180	;
						10'd317	:	dt	<=	186	;
						10'd318	:	dt	<=	192	;
						10'd319	:	dt	<=	197	;
						10'd320	:	dt	<=	201	;
						10'd321	:	dt	<=	203	;
						10'd322	:	dt	<=	207	;
						10'd323	:	dt	<=	208	;
						10'd324	:	dt	<=	210	;
						10'd325	:	dt	<=	255	;
						10'd326	:	dt	<=	255	;
						10'd327	:	dt	<=	204	;
						10'd328	:	dt	<=	216	;
						10'd329	:	dt	<=	206	;
						10'd330	:	dt	<=	200	;
						10'd331	:	dt	<=	216	;
						10'd332	:	dt	<=	213	;
						10'd333	:	dt	<=	213	;
						10'd334	:	dt	<=	212	;
						10'd335	:	dt	<=	211	;
						10'd336	:	dt	<=	121	;
						10'd337	:	dt	<=	124	;
						10'd338	:	dt	<=	132	;
						10'd339	:	dt	<=	145	;
						10'd340	:	dt	<=	157	;
						10'd341	:	dt	<=	167	;
						10'd342	:	dt	<=	174	;
						10'd343	:	dt	<=	176	;
						10'd344	:	dt	<=	181	;
						10'd345	:	dt	<=	188	;
						10'd346	:	dt	<=	193	;
						10'd347	:	dt	<=	199	;
						10'd348	:	dt	<=	204	;
						10'd349	:	dt	<=	202	;
						10'd350	:	dt	<=	206	;
						10'd351	:	dt	<=	207	;
						10'd352	:	dt	<=	232	;
						10'd353	:	dt	<=	255	;
						10'd354	:	dt	<=	255	;
						10'd355	:	dt	<=	255	;
						10'd356	:	dt	<=	255	;
						10'd357	:	dt	<=	175	;
						10'd358	:	dt	<=	165	;
						10'd359	:	dt	<=	227	;
						10'd360	:	dt	<=	213	;
						10'd361	:	dt	<=	215	;
						10'd362	:	dt	<=	214	;
						10'd363	:	dt	<=	213	;
						10'd364	:	dt	<=	121	;
						10'd365	:	dt	<=	125	;
						10'd366	:	dt	<=	133	;
						10'd367	:	dt	<=	146	;
						10'd368	:	dt	<=	157	;
						10'd369	:	dt	<=	169	;
						10'd370	:	dt	<=	175	;
						10'd371	:	dt	<=	177	;
						10'd372	:	dt	<=	183	;
						10'd373	:	dt	<=	189	;
						10'd374	:	dt	<=	194	;
						10'd375	:	dt	<=	202	;
						10'd376	:	dt	<=	200	;
						10'd377	:	dt	<=	215	;
						10'd378	:	dt	<=	236	;
						10'd379	:	dt	<=	244	;
						10'd380	:	dt	<=	255	;
						10'd381	:	dt	<=	218	;
						10'd382	:	dt	<=	241	;
						10'd383	:	dt	<=	230	;
						10'd384	:	dt	<=	218	;
						10'd385	:	dt	<=	158	;
						10'd386	:	dt	<=	135	;
						10'd387	:	dt	<=	201	;
						10'd388	:	dt	<=	214	;
						10'd389	:	dt	<=	217	;
						10'd390	:	dt	<=	216	;
						10'd391	:	dt	<=	215	;
						10'd392	:	dt	<=	122	;
						10'd393	:	dt	<=	126	;
						10'd394	:	dt	<=	135	;
						10'd395	:	dt	<=	147	;
						10'd396	:	dt	<=	159	;
						10'd397	:	dt	<=	170	;
						10'd398	:	dt	<=	177	;
						10'd399	:	dt	<=	180	;
						10'd400	:	dt	<=	185	;
						10'd401	:	dt	<=	190	;
						10'd402	:	dt	<=	197	;
						10'd403	:	dt	<=	198	;
						10'd404	:	dt	<=	218	;
						10'd405	:	dt	<=	251	;
						10'd406	:	dt	<=	244	;
						10'd407	:	dt	<=	251	;
						10'd408	:	dt	<=	255	;
						10'd409	:	dt	<=	227	;
						10'd410	:	dt	<=	254	;
						10'd411	:	dt	<=	255	;
						10'd412	:	dt	<=	226	;
						10'd413	:	dt	<=	155	;
						10'd414	:	dt	<=	122	;
						10'd415	:	dt	<=	172	;
						10'd416	:	dt	<=	196	;
						10'd417	:	dt	<=	224	;
						10'd418	:	dt	<=	216	;
						10'd419	:	dt	<=	217	;
						10'd420	:	dt	<=	122	;
						10'd421	:	dt	<=	125	;
						10'd422	:	dt	<=	135	;
						10'd423	:	dt	<=	148	;
						10'd424	:	dt	<=	160	;
						10'd425	:	dt	<=	171	;
						10'd426	:	dt	<=	178	;
						10'd427	:	dt	<=	181	;
						10'd428	:	dt	<=	186	;
						10'd429	:	dt	<=	193	;
						10'd430	:	dt	<=	196	;
						10'd431	:	dt	<=	209	;
						10'd432	:	dt	<=	251	;
						10'd433	:	dt	<=	232	;
						10'd434	:	dt	<=	224	;
						10'd435	:	dt	<=	230	;
						10'd436	:	dt	<=	230	;
						10'd437	:	dt	<=	211	;
						10'd438	:	dt	<=	232	;
						10'd439	:	dt	<=	246	;
						10'd440	:	dt	<=	210	;
						10'd441	:	dt	<=	144	;
						10'd442	:	dt	<=	114	;
						10'd443	:	dt	<=	138	;
						10'd444	:	dt	<=	153	;
						10'd445	:	dt	<=	229	;
						10'd446	:	dt	<=	219	;
						10'd447	:	dt	<=	218	;
						10'd448	:	dt	<=	123	;
						10'd449	:	dt	<=	125	;
						10'd450	:	dt	<=	134	;
						10'd451	:	dt	<=	148	;
						10'd452	:	dt	<=	161	;
						10'd453	:	dt	<=	172	;
						10'd454	:	dt	<=	180	;
						10'd455	:	dt	<=	181	;
						10'd456	:	dt	<=	186	;
						10'd457	:	dt	<=	195	;
						10'd458	:	dt	<=	193	;
						10'd459	:	dt	<=	255	;
						10'd460	:	dt	<=	255	;
						10'd461	:	dt	<=	249	;
						10'd462	:	dt	<=	239	;
						10'd463	:	dt	<=	240	;
						10'd464	:	dt	<=	228	;
						10'd465	:	dt	<=	215	;
						10'd466	:	dt	<=	215	;
						10'd467	:	dt	<=	180	;
						10'd468	:	dt	<=	163	;
						10'd469	:	dt	<=	144	;
						10'd470	:	dt	<=	109	;
						10'd471	:	dt	<=	141	;
						10'd472	:	dt	<=	124	;
						10'd473	:	dt	<=	174	;
						10'd474	:	dt	<=	226	;
						10'd475	:	dt	<=	220	;
						10'd476	:	dt	<=	123	;
						10'd477	:	dt	<=	125	;
						10'd478	:	dt	<=	135	;
						10'd479	:	dt	<=	148	;
						10'd480	:	dt	<=	161	;
						10'd481	:	dt	<=	172	;
						10'd482	:	dt	<=	180	;
						10'd483	:	dt	<=	182	;
						10'd484	:	dt	<=	187	;
						10'd485	:	dt	<=	195	;
						10'd486	:	dt	<=	199	;
						10'd487	:	dt	<=	255	;
						10'd488	:	dt	<=	255	;
						10'd489	:	dt	<=	251	;
						10'd490	:	dt	<=	215	;
						10'd491	:	dt	<=	216	;
						10'd492	:	dt	<=	231	;
						10'd493	:	dt	<=	227	;
						10'd494	:	dt	<=	216	;
						10'd495	:	dt	<=	164	;
						10'd496	:	dt	<=	141	;
						10'd497	:	dt	<=	152	;
						10'd498	:	dt	<=	100	;
						10'd499	:	dt	<=	138	;
						10'd500	:	dt	<=	141	;
						10'd501	:	dt	<=	132	;
						10'd502	:	dt	<=	205	;
						10'd503	:	dt	<=	226	;
						10'd504	:	dt	<=	122	;
						10'd505	:	dt	<=	124	;
						10'd506	:	dt	<=	135	;
						10'd507	:	dt	<=	150	;
						10'd508	:	dt	<=	161	;
						10'd509	:	dt	<=	173	;
						10'd510	:	dt	<=	180	;
						10'd511	:	dt	<=	182	;
						10'd512	:	dt	<=	187	;
						10'd513	:	dt	<=	194	;
						10'd514	:	dt	<=	202	;
						10'd515	:	dt	<=	255	;
						10'd516	:	dt	<=	255	;
						10'd517	:	dt	<=	236	;
						10'd518	:	dt	<=	189	;
						10'd519	:	dt	<=	160	;
						10'd520	:	dt	<=	172	;
						10'd521	:	dt	<=	191	;
						10'd522	:	dt	<=	195	;
						10'd523	:	dt	<=	150	;
						10'd524	:	dt	<=	148	;
						10'd525	:	dt	<=	149	;
						10'd526	:	dt	<=	93	;
						10'd527	:	dt	<=	134	;
						10'd528	:	dt	<=	143	;
						10'd529	:	dt	<=	150	;
						10'd530	:	dt	<=	217	;
						10'd531	:	dt	<=	224	;
						10'd532	:	dt	<=	122	;
						10'd533	:	dt	<=	125	;
						10'd534	:	dt	<=	136	;
						10'd535	:	dt	<=	150	;
						10'd536	:	dt	<=	162	;
						10'd537	:	dt	<=	175	;
						10'd538	:	dt	<=	180	;
						10'd539	:	dt	<=	182	;
						10'd540	:	dt	<=	187	;
						10'd541	:	dt	<=	194	;
						10'd542	:	dt	<=	205	;
						10'd543	:	dt	<=	255	;
						10'd544	:	dt	<=	255	;
						10'd545	:	dt	<=	206	;
						10'd546	:	dt	<=	154	;
						10'd547	:	dt	<=	133	;
						10'd548	:	dt	<=	104	;
						10'd549	:	dt	<=	201	;
						10'd550	:	dt	<=	194	;
						10'd551	:	dt	<=	141	;
						10'd552	:	dt	<=	156	;
						10'd553	:	dt	<=	127	;
						10'd554	:	dt	<=	112	;
						10'd555	:	dt	<=	146	;
						10'd556	:	dt	<=	141	;
						10'd557	:	dt	<=	183	;
						10'd558	:	dt	<=	231	;
						10'd559	:	dt	<=	223	;
						10'd560	:	dt	<=	122	;
						10'd561	:	dt	<=	124	;
						10'd562	:	dt	<=	138	;
						10'd563	:	dt	<=	151	;
						10'd564	:	dt	<=	162	;
						10'd565	:	dt	<=	174	;
						10'd566	:	dt	<=	181	;
						10'd567	:	dt	<=	184	;
						10'd568	:	dt	<=	191	;
						10'd569	:	dt	<=	194	;
						10'd570	:	dt	<=	208	;
						10'd571	:	dt	<=	255	;
						10'd572	:	dt	<=	255	;
						10'd573	:	dt	<=	201	;
						10'd574	:	dt	<=	157	;
						10'd575	:	dt	<=	119	;
						10'd576	:	dt	<=	127	;
						10'd577	:	dt	<=	202	;
						10'd578	:	dt	<=	171	;
						10'd579	:	dt	<=	144	;
						10'd580	:	dt	<=	132	;
						10'd581	:	dt	<=	98	;
						10'd582	:	dt	<=	130	;
						10'd583	:	dt	<=	153	;
						10'd584	:	dt	<=	155	;
						10'd585	:	dt	<=	224	;
						10'd586	:	dt	<=	228	;
						10'd587	:	dt	<=	228	;
						10'd588	:	dt	<=	121	;
						10'd589	:	dt	<=	124	;
						10'd590	:	dt	<=	137	;
						10'd591	:	dt	<=	151	;
						10'd592	:	dt	<=	163	;
						10'd593	:	dt	<=	176	;
						10'd594	:	dt	<=	182	;
						10'd595	:	dt	<=	184	;
						10'd596	:	dt	<=	192	;
						10'd597	:	dt	<=	193	;
						10'd598	:	dt	<=	217	;
						10'd599	:	dt	<=	255	;
						10'd600	:	dt	<=	250	;
						10'd601	:	dt	<=	198	;
						10'd602	:	dt	<=	162	;
						10'd603	:	dt	<=	129	;
						10'd604	:	dt	<=	119	;
						10'd605	:	dt	<=	130	;
						10'd606	:	dt	<=	131	;
						10'd607	:	dt	<=	113	;
						10'd608	:	dt	<=	105	;
						10'd609	:	dt	<=	114	;
						10'd610	:	dt	<=	131	;
						10'd611	:	dt	<=	143	;
						10'd612	:	dt	<=	187	;
						10'd613	:	dt	<=	237	;
						10'd614	:	dt	<=	228	;
						10'd615	:	dt	<=	229	;
						10'd616	:	dt	<=	119	;
						10'd617	:	dt	<=	122	;
						10'd618	:	dt	<=	136	;
						10'd619	:	dt	<=	151	;
						10'd620	:	dt	<=	162	;
						10'd621	:	dt	<=	174	;
						10'd622	:	dt	<=	180	;
						10'd623	:	dt	<=	182	;
						10'd624	:	dt	<=	190	;
						10'd625	:	dt	<=	191	;
						10'd626	:	dt	<=	225	;
						10'd627	:	dt	<=	255	;
						10'd628	:	dt	<=	244	;
						10'd629	:	dt	<=	196	;
						10'd630	:	dt	<=	162	;
						10'd631	:	dt	<=	126	;
						10'd632	:	dt	<=	94	;
						10'd633	:	dt	<=	100	;
						10'd634	:	dt	<=	106	;
						10'd635	:	dt	<=	118	;
						10'd636	:	dt	<=	136	;
						10'd637	:	dt	<=	137	;
						10'd638	:	dt	<=	136	;
						10'd639	:	dt	<=	142	;
						10'd640	:	dt	<=	217	;
						10'd641	:	dt	<=	232	;
						10'd642	:	dt	<=	229	;
						10'd643	:	dt	<=	229	;
						10'd644	:	dt	<=	118	;
						10'd645	:	dt	<=	121	;
						10'd646	:	dt	<=	135	;
						10'd647	:	dt	<=	149	;
						10'd648	:	dt	<=	163	;
						10'd649	:	dt	<=	174	;
						10'd650	:	dt	<=	182	;
						10'd651	:	dt	<=	183	;
						10'd652	:	dt	<=	192	;
						10'd653	:	dt	<=	192	;
						10'd654	:	dt	<=	236	;
						10'd655	:	dt	<=	255	;
						10'd656	:	dt	<=	238	;
						10'd657	:	dt	<=	198	;
						10'd658	:	dt	<=	162	;
						10'd659	:	dt	<=	135	;
						10'd660	:	dt	<=	113	;
						10'd661	:	dt	<=	126	;
						10'd662	:	dt	<=	139	;
						10'd663	:	dt	<=	145	;
						10'd664	:	dt	<=	151	;
						10'd665	:	dt	<=	144	;
						10'd666	:	dt	<=	133	;
						10'd667	:	dt	<=	180	;
						10'd668	:	dt	<=	235	;
						10'd669	:	dt	<=	231	;
						10'd670	:	dt	<=	230	;
						10'd671	:	dt	<=	229	;
						10'd672	:	dt	<=	117	;
						10'd673	:	dt	<=	121	;
						10'd674	:	dt	<=	134	;
						10'd675	:	dt	<=	149	;
						10'd676	:	dt	<=	162	;
						10'd677	:	dt	<=	175	;
						10'd678	:	dt	<=	182	;
						10'd679	:	dt	<=	184	;
						10'd680	:	dt	<=	193	;
						10'd681	:	dt	<=	193	;
						10'd682	:	dt	<=	234	;
						10'd683	:	dt	<=	255	;
						10'd684	:	dt	<=	230	;
						10'd685	:	dt	<=	194	;
						10'd686	:	dt	<=	165	;
						10'd687	:	dt	<=	141	;
						10'd688	:	dt	<=	124	;
						10'd689	:	dt	<=	130	;
						10'd690	:	dt	<=	150	;
						10'd691	:	dt	<=	154	;
						10'd692	:	dt	<=	154	;
						10'd693	:	dt	<=	139	;
						10'd694	:	dt	<=	152	;
						10'd695	:	dt	<=	234	;
						10'd696	:	dt	<=	233	;
						10'd697	:	dt	<=	232	;
						10'd698	:	dt	<=	232	;
						10'd699	:	dt	<=	231	;
						10'd700	:	dt	<=	115	;
						10'd701	:	dt	<=	119	;
						10'd702	:	dt	<=	132	;
						10'd703	:	dt	<=	148	;
						10'd704	:	dt	<=	163	;
						10'd705	:	dt	<=	174	;
						10'd706	:	dt	<=	182	;
						10'd707	:	dt	<=	184	;
						10'd708	:	dt	<=	192	;
						10'd709	:	dt	<=	193	;
						10'd710	:	dt	<=	236	;
						10'd711	:	dt	<=	255	;
						10'd712	:	dt	<=	220	;
						10'd713	:	dt	<=	195	;
						10'd714	:	dt	<=	170	;
						10'd715	:	dt	<=	147	;
						10'd716	:	dt	<=	136	;
						10'd717	:	dt	<=	132	;
						10'd718	:	dt	<=	152	;
						10'd719	:	dt	<=	157	;
						10'd720	:	dt	<=	156	;
						10'd721	:	dt	<=	133	;
						10'd722	:	dt	<=	192	;
						10'd723	:	dt	<=	242	;
						10'd724	:	dt	<=	231	;
						10'd725	:	dt	<=	233	;
						10'd726	:	dt	<=	232	;
						10'd727	:	dt	<=	231	;
						10'd728	:	dt	<=	112	;
						10'd729	:	dt	<=	116	;
						10'd730	:	dt	<=	130	;
						10'd731	:	dt	<=	146	;
						10'd732	:	dt	<=	161	;
						10'd733	:	dt	<=	174	;
						10'd734	:	dt	<=	180	;
						10'd735	:	dt	<=	183	;
						10'd736	:	dt	<=	191	;
						10'd737	:	dt	<=	193	;
						10'd738	:	dt	<=	245	;
						10'd739	:	dt	<=	248	;
						10'd740	:	dt	<=	224	;
						10'd741	:	dt	<=	211	;
						10'd742	:	dt	<=	184	;
						10'd743	:	dt	<=	158	;
						10'd744	:	dt	<=	143	;
						10'd745	:	dt	<=	133	;
						10'd746	:	dt	<=	149	;
						10'd747	:	dt	<=	155	;
						10'd748	:	dt	<=	146	;
						10'd749	:	dt	<=	158	;
						10'd750	:	dt	<=	232	;
						10'd751	:	dt	<=	235	;
						10'd752	:	dt	<=	234	;
						10'd753	:	dt	<=	232	;
						10'd754	:	dt	<=	232	;
						10'd755	:	dt	<=	232	;
						10'd756	:	dt	<=	114	;
						10'd757	:	dt	<=	118	;
						10'd758	:	dt	<=	130	;
						10'd759	:	dt	<=	145	;
						10'd760	:	dt	<=	158	;
						10'd761	:	dt	<=	171	;
						10'd762	:	dt	<=	178	;
						10'd763	:	dt	<=	181	;
						10'd764	:	dt	<=	190	;
						10'd765	:	dt	<=	195	;
						10'd766	:	dt	<=	255	;
						10'd767	:	dt	<=	254	;
						10'd768	:	dt	<=	237	;
						10'd769	:	dt	<=	224	;
						10'd770	:	dt	<=	197	;
						10'd771	:	dt	<=	163	;
						10'd772	:	dt	<=	147	;
						10'd773	:	dt	<=	138	;
						10'd774	:	dt	<=	148	;
						10'd775	:	dt	<=	149	;
						10'd776	:	dt	<=	149	;
						10'd777	:	dt	<=	216	;
						10'd778	:	dt	<=	238	;
						10'd779	:	dt	<=	231	;
						10'd780	:	dt	<=	232	;
						10'd781	:	dt	<=	231	;
						10'd782	:	dt	<=	232	;
						10'd783	:	dt	<=	231	;
					endcase
				end
				5'd24	:	begin
					case (cnt)
						10'd0	:	dt	<=	158	;
						10'd1	:	dt	<=	160	;
						10'd2	:	dt	<=	163	;
						10'd3	:	dt	<=	163	;
						10'd4	:	dt	<=	164	;
						10'd5	:	dt	<=	165	;
						10'd6	:	dt	<=	166	;
						10'd7	:	dt	<=	166	;
						10'd8	:	dt	<=	167	;
						10'd9	:	dt	<=	167	;
						10'd10	:	dt	<=	166	;
						10'd11	:	dt	<=	167	;
						10'd12	:	dt	<=	166	;
						10'd13	:	dt	<=	165	;
						10'd14	:	dt	<=	165	;
						10'd15	:	dt	<=	163	;
						10'd16	:	dt	<=	162	;
						10'd17	:	dt	<=	162	;
						10'd18	:	dt	<=	161	;
						10'd19	:	dt	<=	161	;
						10'd20	:	dt	<=	160	;
						10'd21	:	dt	<=	158	;
						10'd22	:	dt	<=	157	;
						10'd23	:	dt	<=	156	;
						10'd24	:	dt	<=	155	;
						10'd25	:	dt	<=	153	;
						10'd26	:	dt	<=	152	;
						10'd27	:	dt	<=	152	;
						10'd28	:	dt	<=	159	;
						10'd29	:	dt	<=	162	;
						10'd30	:	dt	<=	165	;
						10'd31	:	dt	<=	164	;
						10'd32	:	dt	<=	165	;
						10'd33	:	dt	<=	166	;
						10'd34	:	dt	<=	167	;
						10'd35	:	dt	<=	168	;
						10'd36	:	dt	<=	168	;
						10'd37	:	dt	<=	168	;
						10'd38	:	dt	<=	168	;
						10'd39	:	dt	<=	168	;
						10'd40	:	dt	<=	168	;
						10'd41	:	dt	<=	166	;
						10'd42	:	dt	<=	166	;
						10'd43	:	dt	<=	166	;
						10'd44	:	dt	<=	164	;
						10'd45	:	dt	<=	164	;
						10'd46	:	dt	<=	164	;
						10'd47	:	dt	<=	164	;
						10'd48	:	dt	<=	161	;
						10'd49	:	dt	<=	160	;
						10'd50	:	dt	<=	160	;
						10'd51	:	dt	<=	159	;
						10'd52	:	dt	<=	159	;
						10'd53	:	dt	<=	156	;
						10'd54	:	dt	<=	156	;
						10'd55	:	dt	<=	154	;
						10'd56	:	dt	<=	160	;
						10'd57	:	dt	<=	163	;
						10'd58	:	dt	<=	165	;
						10'd59	:	dt	<=	166	;
						10'd60	:	dt	<=	168	;
						10'd61	:	dt	<=	168	;
						10'd62	:	dt	<=	169	;
						10'd63	:	dt	<=	170	;
						10'd64	:	dt	<=	171	;
						10'd65	:	dt	<=	170	;
						10'd66	:	dt	<=	170	;
						10'd67	:	dt	<=	171	;
						10'd68	:	dt	<=	171	;
						10'd69	:	dt	<=	170	;
						10'd70	:	dt	<=	168	;
						10'd71	:	dt	<=	167	;
						10'd72	:	dt	<=	166	;
						10'd73	:	dt	<=	167	;
						10'd74	:	dt	<=	165	;
						10'd75	:	dt	<=	164	;
						10'd76	:	dt	<=	164	;
						10'd77	:	dt	<=	162	;
						10'd78	:	dt	<=	161	;
						10'd79	:	dt	<=	161	;
						10'd80	:	dt	<=	160	;
						10'd81	:	dt	<=	159	;
						10'd82	:	dt	<=	157	;
						10'd83	:	dt	<=	156	;
						10'd84	:	dt	<=	162	;
						10'd85	:	dt	<=	163	;
						10'd86	:	dt	<=	166	;
						10'd87	:	dt	<=	167	;
						10'd88	:	dt	<=	169	;
						10'd89	:	dt	<=	169	;
						10'd90	:	dt	<=	170	;
						10'd91	:	dt	<=	171	;
						10'd92	:	dt	<=	171	;
						10'd93	:	dt	<=	170	;
						10'd94	:	dt	<=	171	;
						10'd95	:	dt	<=	171	;
						10'd96	:	dt	<=	171	;
						10'd97	:	dt	<=	172	;
						10'd98	:	dt	<=	170	;
						10'd99	:	dt	<=	169	;
						10'd100	:	dt	<=	169	;
						10'd101	:	dt	<=	167	;
						10'd102	:	dt	<=	165	;
						10'd103	:	dt	<=	166	;
						10'd104	:	dt	<=	165	;
						10'd105	:	dt	<=	165	;
						10'd106	:	dt	<=	164	;
						10'd107	:	dt	<=	163	;
						10'd108	:	dt	<=	161	;
						10'd109	:	dt	<=	160	;
						10'd110	:	dt	<=	159	;
						10'd111	:	dt	<=	158	;
						10'd112	:	dt	<=	163	;
						10'd113	:	dt	<=	164	;
						10'd114	:	dt	<=	167	;
						10'd115	:	dt	<=	168	;
						10'd116	:	dt	<=	168	;
						10'd117	:	dt	<=	167	;
						10'd118	:	dt	<=	171	;
						10'd119	:	dt	<=	174	;
						10'd120	:	dt	<=	173	;
						10'd121	:	dt	<=	172	;
						10'd122	:	dt	<=	172	;
						10'd123	:	dt	<=	172	;
						10'd124	:	dt	<=	172	;
						10'd125	:	dt	<=	172	;
						10'd126	:	dt	<=	170	;
						10'd127	:	dt	<=	169	;
						10'd128	:	dt	<=	169	;
						10'd129	:	dt	<=	167	;
						10'd130	:	dt	<=	167	;
						10'd131	:	dt	<=	167	;
						10'd132	:	dt	<=	166	;
						10'd133	:	dt	<=	165	;
						10'd134	:	dt	<=	165	;
						10'd135	:	dt	<=	164	;
						10'd136	:	dt	<=	163	;
						10'd137	:	dt	<=	161	;
						10'd138	:	dt	<=	160	;
						10'd139	:	dt	<=	159	;
						10'd140	:	dt	<=	165	;
						10'd141	:	dt	<=	165	;
						10'd142	:	dt	<=	169	;
						10'd143	:	dt	<=	166	;
						10'd144	:	dt	<=	181	;
						10'd145	:	dt	<=	153	;
						10'd146	:	dt	<=	129	;
						10'd147	:	dt	<=	178	;
						10'd148	:	dt	<=	173	;
						10'd149	:	dt	<=	174	;
						10'd150	:	dt	<=	174	;
						10'd151	:	dt	<=	173	;
						10'd152	:	dt	<=	173	;
						10'd153	:	dt	<=	173	;
						10'd154	:	dt	<=	172	;
						10'd155	:	dt	<=	171	;
						10'd156	:	dt	<=	171	;
						10'd157	:	dt	<=	169	;
						10'd158	:	dt	<=	168	;
						10'd159	:	dt	<=	168	;
						10'd160	:	dt	<=	168	;
						10'd161	:	dt	<=	167	;
						10'd162	:	dt	<=	166	;
						10'd163	:	dt	<=	164	;
						10'd164	:	dt	<=	164	;
						10'd165	:	dt	<=	163	;
						10'd166	:	dt	<=	162	;
						10'd167	:	dt	<=	161	;
						10'd168	:	dt	<=	166	;
						10'd169	:	dt	<=	167	;
						10'd170	:	dt	<=	170	;
						10'd171	:	dt	<=	167	;
						10'd172	:	dt	<=	190	;
						10'd173	:	dt	<=	132	;
						10'd174	:	dt	<=	112	;
						10'd175	:	dt	<=	181	;
						10'd176	:	dt	<=	173	;
						10'd177	:	dt	<=	174	;
						10'd178	:	dt	<=	174	;
						10'd179	:	dt	<=	175	;
						10'd180	:	dt	<=	174	;
						10'd181	:	dt	<=	174	;
						10'd182	:	dt	<=	173	;
						10'd183	:	dt	<=	172	;
						10'd184	:	dt	<=	172	;
						10'd185	:	dt	<=	171	;
						10'd186	:	dt	<=	169	;
						10'd187	:	dt	<=	169	;
						10'd188	:	dt	<=	169	;
						10'd189	:	dt	<=	168	;
						10'd190	:	dt	<=	167	;
						10'd191	:	dt	<=	166	;
						10'd192	:	dt	<=	165	;
						10'd193	:	dt	<=	164	;
						10'd194	:	dt	<=	163	;
						10'd195	:	dt	<=	162	;
						10'd196	:	dt	<=	166	;
						10'd197	:	dt	<=	168	;
						10'd198	:	dt	<=	170	;
						10'd199	:	dt	<=	171	;
						10'd200	:	dt	<=	186	;
						10'd201	:	dt	<=	110	;
						10'd202	:	dt	<=	127	;
						10'd203	:	dt	<=	182	;
						10'd204	:	dt	<=	173	;
						10'd205	:	dt	<=	175	;
						10'd206	:	dt	<=	176	;
						10'd207	:	dt	<=	176	;
						10'd208	:	dt	<=	177	;
						10'd209	:	dt	<=	174	;
						10'd210	:	dt	<=	173	;
						10'd211	:	dt	<=	172	;
						10'd212	:	dt	<=	172	;
						10'd213	:	dt	<=	171	;
						10'd214	:	dt	<=	171	;
						10'd215	:	dt	<=	170	;
						10'd216	:	dt	<=	170	;
						10'd217	:	dt	<=	169	;
						10'd218	:	dt	<=	168	;
						10'd219	:	dt	<=	167	;
						10'd220	:	dt	<=	166	;
						10'd221	:	dt	<=	165	;
						10'd222	:	dt	<=	164	;
						10'd223	:	dt	<=	163	;
						10'd224	:	dt	<=	168	;
						10'd225	:	dt	<=	170	;
						10'd226	:	dt	<=	170	;
						10'd227	:	dt	<=	177	;
						10'd228	:	dt	<=	184	;
						10'd229	:	dt	<=	109	;
						10'd230	:	dt	<=	137	;
						10'd231	:	dt	<=	183	;
						10'd232	:	dt	<=	175	;
						10'd233	:	dt	<=	177	;
						10'd234	:	dt	<=	176	;
						10'd235	:	dt	<=	174	;
						10'd236	:	dt	<=	170	;
						10'd237	:	dt	<=	177	;
						10'd238	:	dt	<=	176	;
						10'd239	:	dt	<=	173	;
						10'd240	:	dt	<=	174	;
						10'd241	:	dt	<=	173	;
						10'd242	:	dt	<=	172	;
						10'd243	:	dt	<=	172	;
						10'd244	:	dt	<=	171	;
						10'd245	:	dt	<=	170	;
						10'd246	:	dt	<=	168	;
						10'd247	:	dt	<=	167	;
						10'd248	:	dt	<=	166	;
						10'd249	:	dt	<=	167	;
						10'd250	:	dt	<=	165	;
						10'd251	:	dt	<=	165	;
						10'd252	:	dt	<=	170	;
						10'd253	:	dt	<=	171	;
						10'd254	:	dt	<=	172	;
						10'd255	:	dt	<=	181	;
						10'd256	:	dt	<=	183	;
						10'd257	:	dt	<=	106	;
						10'd258	:	dt	<=	141	;
						10'd259	:	dt	<=	190	;
						10'd260	:	dt	<=	177	;
						10'd261	:	dt	<=	177	;
						10'd262	:	dt	<=	183	;
						10'd263	:	dt	<=	181	;
						10'd264	:	dt	<=	149	;
						10'd265	:	dt	<=	121	;
						10'd266	:	dt	<=	175	;
						10'd267	:	dt	<=	177	;
						10'd268	:	dt	<=	173	;
						10'd269	:	dt	<=	174	;
						10'd270	:	dt	<=	173	;
						10'd271	:	dt	<=	173	;
						10'd272	:	dt	<=	174	;
						10'd273	:	dt	<=	173	;
						10'd274	:	dt	<=	174	;
						10'd275	:	dt	<=	171	;
						10'd276	:	dt	<=	167	;
						10'd277	:	dt	<=	167	;
						10'd278	:	dt	<=	167	;
						10'd279	:	dt	<=	166	;
						10'd280	:	dt	<=	171	;
						10'd281	:	dt	<=	172	;
						10'd282	:	dt	<=	172	;
						10'd283	:	dt	<=	183	;
						10'd284	:	dt	<=	170	;
						10'd285	:	dt	<=	125	;
						10'd286	:	dt	<=	146	;
						10'd287	:	dt	<=	158	;
						10'd288	:	dt	<=	181	;
						10'd289	:	dt	<=	144	;
						10'd290	:	dt	<=	144	;
						10'd291	:	dt	<=	183	;
						10'd292	:	dt	<=	166	;
						10'd293	:	dt	<=	119	;
						10'd294	:	dt	<=	102	;
						10'd295	:	dt	<=	176	;
						10'd296	:	dt	<=	177	;
						10'd297	:	dt	<=	175	;
						10'd298	:	dt	<=	175	;
						10'd299	:	dt	<=	173	;
						10'd300	:	dt	<=	164	;
						10'd301	:	dt	<=	151	;
						10'd302	:	dt	<=	143	;
						10'd303	:	dt	<=	164	;
						10'd304	:	dt	<=	172	;
						10'd305	:	dt	<=	168	;
						10'd306	:	dt	<=	168	;
						10'd307	:	dt	<=	167	;
						10'd308	:	dt	<=	170	;
						10'd309	:	dt	<=	175	;
						10'd310	:	dt	<=	173	;
						10'd311	:	dt	<=	186	;
						10'd312	:	dt	<=	180	;
						10'd313	:	dt	<=	185	;
						10'd314	:	dt	<=	179	;
						10'd315	:	dt	<=	150	;
						10'd316	:	dt	<=	196	;
						10'd317	:	dt	<=	149	;
						10'd318	:	dt	<=	105	;
						10'd319	:	dt	<=	172	;
						10'd320	:	dt	<=	177	;
						10'd321	:	dt	<=	131	;
						10'd322	:	dt	<=	68	;
						10'd323	:	dt	<=	124	;
						10'd324	:	dt	<=	184	;
						10'd325	:	dt	<=	175	;
						10'd326	:	dt	<=	172	;
						10'd327	:	dt	<=	153	;
						10'd328	:	dt	<=	116	;
						10'd329	:	dt	<=	101	;
						10'd330	:	dt	<=	86	;
						10'd331	:	dt	<=	117	;
						10'd332	:	dt	<=	178	;
						10'd333	:	dt	<=	170	;
						10'd334	:	dt	<=	170	;
						10'd335	:	dt	<=	167	;
						10'd336	:	dt	<=	171	;
						10'd337	:	dt	<=	176	;
						10'd338	:	dt	<=	175	;
						10'd339	:	dt	<=	185	;
						10'd340	:	dt	<=	184	;
						10'd341	:	dt	<=	205	;
						10'd342	:	dt	<=	180	;
						10'd343	:	dt	<=	172	;
						10'd344	:	dt	<=	196	;
						10'd345	:	dt	<=	164	;
						10'd346	:	dt	<=	101	;
						10'd347	:	dt	<=	165	;
						10'd348	:	dt	<=	171	;
						10'd349	:	dt	<=	120	;
						10'd350	:	dt	<=	69	;
						10'd351	:	dt	<=	89	;
						10'd352	:	dt	<=	177	;
						10'd353	:	dt	<=	174	;
						10'd354	:	dt	<=	166	;
						10'd355	:	dt	<=	126	;
						10'd356	:	dt	<=	88	;
						10'd357	:	dt	<=	90	;
						10'd358	:	dt	<=	116	;
						10'd359	:	dt	<=	145	;
						10'd360	:	dt	<=	173	;
						10'd361	:	dt	<=	171	;
						10'd362	:	dt	<=	170	;
						10'd363	:	dt	<=	168	;
						10'd364	:	dt	<=	174	;
						10'd365	:	dt	<=	176	;
						10'd366	:	dt	<=	176	;
						10'd367	:	dt	<=	187	;
						10'd368	:	dt	<=	179	;
						10'd369	:	dt	<=	212	;
						10'd370	:	dt	<=	185	;
						10'd371	:	dt	<=	183	;
						10'd372	:	dt	<=	203	;
						10'd373	:	dt	<=	158	;
						10'd374	:	dt	<=	86	;
						10'd375	:	dt	<=	127	;
						10'd376	:	dt	<=	136	;
						10'd377	:	dt	<=	95	;
						10'd378	:	dt	<=	52	;
						10'd379	:	dt	<=	64	;
						10'd380	:	dt	<=	155	;
						10'd381	:	dt	<=	175	;
						10'd382	:	dt	<=	149	;
						10'd383	:	dt	<=	104	;
						10'd384	:	dt	<=	86	;
						10'd385	:	dt	<=	156	;
						10'd386	:	dt	<=	178	;
						10'd387	:	dt	<=	175	;
						10'd388	:	dt	<=	172	;
						10'd389	:	dt	<=	172	;
						10'd390	:	dt	<=	171	;
						10'd391	:	dt	<=	170	;
						10'd392	:	dt	<=	175	;
						10'd393	:	dt	<=	179	;
						10'd394	:	dt	<=	176	;
						10'd395	:	dt	<=	191	;
						10'd396	:	dt	<=	207	;
						10'd397	:	dt	<=	209	;
						10'd398	:	dt	<=	177	;
						10'd399	:	dt	<=	186	;
						10'd400	:	dt	<=	211	;
						10'd401	:	dt	<=	146	;
						10'd402	:	dt	<=	92	;
						10'd403	:	dt	<=	40	;
						10'd404	:	dt	<=	91	;
						10'd405	:	dt	<=	126	;
						10'd406	:	dt	<=	100	;
						10'd407	:	dt	<=	110	;
						10'd408	:	dt	<=	152	;
						10'd409	:	dt	<=	152	;
						10'd410	:	dt	<=	117	;
						10'd411	:	dt	<=	88	;
						10'd412	:	dt	<=	142	;
						10'd413	:	dt	<=	186	;
						10'd414	:	dt	<=	174	;
						10'd415	:	dt	<=	175	;
						10'd416	:	dt	<=	174	;
						10'd417	:	dt	<=	173	;
						10'd418	:	dt	<=	172	;
						10'd419	:	dt	<=	171	;
						10'd420	:	dt	<=	175	;
						10'd421	:	dt	<=	179	;
						10'd422	:	dt	<=	178	;
						10'd423	:	dt	<=	196	;
						10'd424	:	dt	<=	202	;
						10'd425	:	dt	<=	190	;
						10'd426	:	dt	<=	157	;
						10'd427	:	dt	<=	144	;
						10'd428	:	dt	<=	177	;
						10'd429	:	dt	<=	119	;
						10'd430	:	dt	<=	76	;
						10'd431	:	dt	<=	73	;
						10'd432	:	dt	<=	161	;
						10'd433	:	dt	<=	179	;
						10'd434	:	dt	<=	165	;
						10'd435	:	dt	<=	154	;
						10'd436	:	dt	<=	150	;
						10'd437	:	dt	<=	122	;
						10'd438	:	dt	<=	87	;
						10'd439	:	dt	<=	113	;
						10'd440	:	dt	<=	183	;
						10'd441	:	dt	<=	177	;
						10'd442	:	dt	<=	179	;
						10'd443	:	dt	<=	177	;
						10'd444	:	dt	<=	176	;
						10'd445	:	dt	<=	175	;
						10'd446	:	dt	<=	173	;
						10'd447	:	dt	<=	172	;
						10'd448	:	dt	<=	176	;
						10'd449	:	dt	<=	178	;
						10'd450	:	dt	<=	184	;
						10'd451	:	dt	<=	194	;
						10'd452	:	dt	<=	169	;
						10'd453	:	dt	<=	172	;
						10'd454	:	dt	<=	147	;
						10'd455	:	dt	<=	107	;
						10'd456	:	dt	<=	103	;
						10'd457	:	dt	<=	107	;
						10'd458	:	dt	<=	151	;
						10'd459	:	dt	<=	198	;
						10'd460	:	dt	<=	193	;
						10'd461	:	dt	<=	174	;
						10'd462	:	dt	<=	159	;
						10'd463	:	dt	<=	140	;
						10'd464	:	dt	<=	130	;
						10'd465	:	dt	<=	113	;
						10'd466	:	dt	<=	88	;
						10'd467	:	dt	<=	168	;
						10'd468	:	dt	<=	182	;
						10'd469	:	dt	<=	179	;
						10'd470	:	dt	<=	180	;
						10'd471	:	dt	<=	178	;
						10'd472	:	dt	<=	178	;
						10'd473	:	dt	<=	176	;
						10'd474	:	dt	<=	174	;
						10'd475	:	dt	<=	173	;
						10'd476	:	dt	<=	177	;
						10'd477	:	dt	<=	177	;
						10'd478	:	dt	<=	188	;
						10'd479	:	dt	<=	208	;
						10'd480	:	dt	<=	180	;
						10'd481	:	dt	<=	166	;
						10'd482	:	dt	<=	152	;
						10'd483	:	dt	<=	135	;
						10'd484	:	dt	<=	101	;
						10'd485	:	dt	<=	197	;
						10'd486	:	dt	<=	214	;
						10'd487	:	dt	<=	199	;
						10'd488	:	dt	<=	189	;
						10'd489	:	dt	<=	171	;
						10'd490	:	dt	<=	144	;
						10'd491	:	dt	<=	127	;
						10'd492	:	dt	<=	113	;
						10'd493	:	dt	<=	101	;
						10'd494	:	dt	<=	130	;
						10'd495	:	dt	<=	188	;
						10'd496	:	dt	<=	179	;
						10'd497	:	dt	<=	181	;
						10'd498	:	dt	<=	179	;
						10'd499	:	dt	<=	178	;
						10'd500	:	dt	<=	179	;
						10'd501	:	dt	<=	176	;
						10'd502	:	dt	<=	175	;
						10'd503	:	dt	<=	174	;
						10'd504	:	dt	<=	178	;
						10'd505	:	dt	<=	176	;
						10'd506	:	dt	<=	195	;
						10'd507	:	dt	<=	214	;
						10'd508	:	dt	<=	190	;
						10'd509	:	dt	<=	168	;
						10'd510	:	dt	<=	151	;
						10'd511	:	dt	<=	161	;
						10'd512	:	dt	<=	203	;
						10'd513	:	dt	<=	220	;
						10'd514	:	dt	<=	201	;
						10'd515	:	dt	<=	195	;
						10'd516	:	dt	<=	184	;
						10'd517	:	dt	<=	159	;
						10'd518	:	dt	<=	132	;
						10'd519	:	dt	<=	111	;
						10'd520	:	dt	<=	108	;
						10'd521	:	dt	<=	101	;
						10'd522	:	dt	<=	176	;
						10'd523	:	dt	<=	186	;
						10'd524	:	dt	<=	182	;
						10'd525	:	dt	<=	181	;
						10'd526	:	dt	<=	180	;
						10'd527	:	dt	<=	179	;
						10'd528	:	dt	<=	179	;
						10'd529	:	dt	<=	177	;
						10'd530	:	dt	<=	175	;
						10'd531	:	dt	<=	176	;
						10'd532	:	dt	<=	179	;
						10'd533	:	dt	<=	177	;
						10'd534	:	dt	<=	204	;
						10'd535	:	dt	<=	218	;
						10'd536	:	dt	<=	195	;
						10'd537	:	dt	<=	182	;
						10'd538	:	dt	<=	182	;
						10'd539	:	dt	<=	209	;
						10'd540	:	dt	<=	221	;
						10'd541	:	dt	<=	212	;
						10'd542	:	dt	<=	204	;
						10'd543	:	dt	<=	190	;
						10'd544	:	dt	<=	171	;
						10'd545	:	dt	<=	144	;
						10'd546	:	dt	<=	114	;
						10'd547	:	dt	<=	110	;
						10'd548	:	dt	<=	92	;
						10'd549	:	dt	<=	129	;
						10'd550	:	dt	<=	192	;
						10'd551	:	dt	<=	184	;
						10'd552	:	dt	<=	185	;
						10'd553	:	dt	<=	182	;
						10'd554	:	dt	<=	181	;
						10'd555	:	dt	<=	180	;
						10'd556	:	dt	<=	180	;
						10'd557	:	dt	<=	178	;
						10'd558	:	dt	<=	178	;
						10'd559	:	dt	<=	177	;
						10'd560	:	dt	<=	180	;
						10'd561	:	dt	<=	177	;
						10'd562	:	dt	<=	209	;
						10'd563	:	dt	<=	219	;
						10'd564	:	dt	<=	200	;
						10'd565	:	dt	<=	190	;
						10'd566	:	dt	<=	206	;
						10'd567	:	dt	<=	221	;
						10'd568	:	dt	<=	220	;
						10'd569	:	dt	<=	208	;
						10'd570	:	dt	<=	200	;
						10'd571	:	dt	<=	178	;
						10'd572	:	dt	<=	153	;
						10'd573	:	dt	<=	124	;
						10'd574	:	dt	<=	110	;
						10'd575	:	dt	<=	100	;
						10'd576	:	dt	<=	100	;
						10'd577	:	dt	<=	181	;
						10'd578	:	dt	<=	187	;
						10'd579	:	dt	<=	185	;
						10'd580	:	dt	<=	186	;
						10'd581	:	dt	<=	183	;
						10'd582	:	dt	<=	182	;
						10'd583	:	dt	<=	181	;
						10'd584	:	dt	<=	180	;
						10'd585	:	dt	<=	181	;
						10'd586	:	dt	<=	179	;
						10'd587	:	dt	<=	178	;
						10'd588	:	dt	<=	182	;
						10'd589	:	dt	<=	178	;
						10'd590	:	dt	<=	209	;
						10'd591	:	dt	<=	225	;
						10'd592	:	dt	<=	204	;
						10'd593	:	dt	<=	192	;
						10'd594	:	dt	<=	211	;
						10'd595	:	dt	<=	218	;
						10'd596	:	dt	<=	204	;
						10'd597	:	dt	<=	186	;
						10'd598	:	dt	<=	179	;
						10'd599	:	dt	<=	159	;
						10'd600	:	dt	<=	131	;
						10'd601	:	dt	<=	114	;
						10'd602	:	dt	<=	102	;
						10'd603	:	dt	<=	96	;
						10'd604	:	dt	<=	169	;
						10'd605	:	dt	<=	192	;
						10'd606	:	dt	<=	187	;
						10'd607	:	dt	<=	187	;
						10'd608	:	dt	<=	186	;
						10'd609	:	dt	<=	185	;
						10'd610	:	dt	<=	184	;
						10'd611	:	dt	<=	183	;
						10'd612	:	dt	<=	181	;
						10'd613	:	dt	<=	181	;
						10'd614	:	dt	<=	180	;
						10'd615	:	dt	<=	178	;
						10'd616	:	dt	<=	181	;
						10'd617	:	dt	<=	178	;
						10'd618	:	dt	<=	203	;
						10'd619	:	dt	<=	228	;
						10'd620	:	dt	<=	208	;
						10'd621	:	dt	<=	190	;
						10'd622	:	dt	<=	200	;
						10'd623	:	dt	<=	203	;
						10'd624	:	dt	<=	194	;
						10'd625	:	dt	<=	169	;
						10'd626	:	dt	<=	157	;
						10'd627	:	dt	<=	138	;
						10'd628	:	dt	<=	116	;
						10'd629	:	dt	<=	105	;
						10'd630	:	dt	<=	100	;
						10'd631	:	dt	<=	169	;
						10'd632	:	dt	<=	195	;
						10'd633	:	dt	<=	188	;
						10'd634	:	dt	<=	189	;
						10'd635	:	dt	<=	187	;
						10'd636	:	dt	<=	186	;
						10'd637	:	dt	<=	186	;
						10'd638	:	dt	<=	184	;
						10'd639	:	dt	<=	184	;
						10'd640	:	dt	<=	182	;
						10'd641	:	dt	<=	181	;
						10'd642	:	dt	<=	180	;
						10'd643	:	dt	<=	179	;
						10'd644	:	dt	<=	182	;
						10'd645	:	dt	<=	182	;
						10'd646	:	dt	<=	195	;
						10'd647	:	dt	<=	210	;
						10'd648	:	dt	<=	194	;
						10'd649	:	dt	<=	189	;
						10'd650	:	dt	<=	204	;
						10'd651	:	dt	<=	206	;
						10'd652	:	dt	<=	194	;
						10'd653	:	dt	<=	171	;
						10'd654	:	dt	<=	155	;
						10'd655	:	dt	<=	129	;
						10'd656	:	dt	<=	105	;
						10'd657	:	dt	<=	83	;
						10'd658	:	dt	<=	159	;
						10'd659	:	dt	<=	199	;
						10'd660	:	dt	<=	191	;
						10'd661	:	dt	<=	191	;
						10'd662	:	dt	<=	189	;
						10'd663	:	dt	<=	188	;
						10'd664	:	dt	<=	188	;
						10'd665	:	dt	<=	187	;
						10'd666	:	dt	<=	186	;
						10'd667	:	dt	<=	185	;
						10'd668	:	dt	<=	183	;
						10'd669	:	dt	<=	183	;
						10'd670	:	dt	<=	181	;
						10'd671	:	dt	<=	180	;
						10'd672	:	dt	<=	182	;
						10'd673	:	dt	<=	184	;
						10'd674	:	dt	<=	188	;
						10'd675	:	dt	<=	195	;
						10'd676	:	dt	<=	188	;
						10'd677	:	dt	<=	197	;
						10'd678	:	dt	<=	202	;
						10'd679	:	dt	<=	194	;
						10'd680	:	dt	<=	190	;
						10'd681	:	dt	<=	163	;
						10'd682	:	dt	<=	143	;
						10'd683	:	dt	<=	118	;
						10'd684	:	dt	<=	78	;
						10'd685	:	dt	<=	108	;
						10'd686	:	dt	<=	198	;
						10'd687	:	dt	<=	192	;
						10'd688	:	dt	<=	193	;
						10'd689	:	dt	<=	191	;
						10'd690	:	dt	<=	191	;
						10'd691	:	dt	<=	189	;
						10'd692	:	dt	<=	189	;
						10'd693	:	dt	<=	188	;
						10'd694	:	dt	<=	187	;
						10'd695	:	dt	<=	185	;
						10'd696	:	dt	<=	184	;
						10'd697	:	dt	<=	184	;
						10'd698	:	dt	<=	181	;
						10'd699	:	dt	<=	180	;
						10'd700	:	dt	<=	182	;
						10'd701	:	dt	<=	185	;
						10'd702	:	dt	<=	187	;
						10'd703	:	dt	<=	201	;
						10'd704	:	dt	<=	210	;
						10'd705	:	dt	<=	201	;
						10'd706	:	dt	<=	196	;
						10'd707	:	dt	<=	184	;
						10'd708	:	dt	<=	186	;
						10'd709	:	dt	<=	159	;
						10'd710	:	dt	<=	134	;
						10'd711	:	dt	<=	104	;
						10'd712	:	dt	<=	69	;
						10'd713	:	dt	<=	155	;
						10'd714	:	dt	<=	200	;
						10'd715	:	dt	<=	193	;
						10'd716	:	dt	<=	194	;
						10'd717	:	dt	<=	193	;
						10'd718	:	dt	<=	193	;
						10'd719	:	dt	<=	190	;
						10'd720	:	dt	<=	189	;
						10'd721	:	dt	<=	188	;
						10'd722	:	dt	<=	187	;
						10'd723	:	dt	<=	187	;
						10'd724	:	dt	<=	185	;
						10'd725	:	dt	<=	183	;
						10'd726	:	dt	<=	183	;
						10'd727	:	dt	<=	182	;
						10'd728	:	dt	<=	182	;
						10'd729	:	dt	<=	184	;
						10'd730	:	dt	<=	186	;
						10'd731	:	dt	<=	213	;
						10'd732	:	dt	<=	212	;
						10'd733	:	dt	<=	187	;
						10'd734	:	dt	<=	194	;
						10'd735	:	dt	<=	183	;
						10'd736	:	dt	<=	173	;
						10'd737	:	dt	<=	153	;
						10'd738	:	dt	<=	132	;
						10'd739	:	dt	<=	93	;
						10'd740	:	dt	<=	80	;
						10'd741	:	dt	<=	183	;
						10'd742	:	dt	<=	198	;
						10'd743	:	dt	<=	195	;
						10'd744	:	dt	<=	194	;
						10'd745	:	dt	<=	195	;
						10'd746	:	dt	<=	194	;
						10'd747	:	dt	<=	191	;
						10'd748	:	dt	<=	190	;
						10'd749	:	dt	<=	189	;
						10'd750	:	dt	<=	188	;
						10'd751	:	dt	<=	187	;
						10'd752	:	dt	<=	186	;
						10'd753	:	dt	<=	186	;
						10'd754	:	dt	<=	184	;
						10'd755	:	dt	<=	181	;
						10'd756	:	dt	<=	180	;
						10'd757	:	dt	<=	183	;
						10'd758	:	dt	<=	185	;
						10'd759	:	dt	<=	220	;
						10'd760	:	dt	<=	210	;
						10'd761	:	dt	<=	177	;
						10'd762	:	dt	<=	200	;
						10'd763	:	dt	<=	178	;
						10'd764	:	dt	<=	162	;
						10'd765	:	dt	<=	153	;
						10'd766	:	dt	<=	125	;
						10'd767	:	dt	<=	96	;
						10'd768	:	dt	<=	83	;
						10'd769	:	dt	<=	186	;
						10'd770	:	dt	<=	196	;
						10'd771	:	dt	<=	193	;
						10'd772	:	dt	<=	193	;
						10'd773	:	dt	<=	194	;
						10'd774	:	dt	<=	192	;
						10'd775	:	dt	<=	191	;
						10'd776	:	dt	<=	189	;
						10'd777	:	dt	<=	188	;
						10'd778	:	dt	<=	188	;
						10'd779	:	dt	<=	187	;
						10'd780	:	dt	<=	186	;
						10'd781	:	dt	<=	185	;
						10'd782	:	dt	<=	183	;
						10'd783	:	dt	<=	182	;
					endcase
				end
			endcase
		end
	end

	assign	q_data = dt;
	
endmodule
